magic
tech sky130A
magscale 1 2
timestamp 1677819468
<< viali >>
rect 5181 8041 5215 8075
rect 5917 8041 5951 8075
rect 3985 7837 4019 7871
rect 4997 7837 5031 7871
rect 5733 7837 5767 7871
rect 3341 7769 3375 7803
rect 2053 7701 2087 7735
rect 4169 7701 4203 7735
rect 1685 7497 1719 7531
rect 1869 7361 1903 7395
rect 2329 7361 2363 7395
rect 2973 7361 3007 7395
rect 2421 7157 2455 7191
rect 4261 7157 4295 7191
rect 2053 6817 2087 6851
rect 4261 6749 4295 6783
rect 4445 6749 4479 6783
rect 5181 6749 5215 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 6561 6749 6595 6783
rect 2320 6681 2354 6715
rect 3433 6613 3467 6647
rect 4077 6613 4111 6647
rect 4997 6613 5031 6647
rect 5733 6613 5767 6647
rect 6377 6613 6411 6647
rect 4629 6409 4663 6443
rect 3166 6273 3200 6307
rect 3433 6273 3467 6307
rect 3893 6273 3927 6307
rect 5742 6273 5776 6307
rect 6009 6205 6043 6239
rect 2053 6069 2087 6103
rect 3985 6069 4019 6103
rect 5273 5865 5307 5899
rect 3433 5729 3467 5763
rect 4813 5729 4847 5763
rect 5733 5729 5767 5763
rect 3985 5661 4019 5695
rect 4721 5661 4755 5695
rect 4997 5661 5031 5695
rect 5089 5661 5123 5695
rect 6009 5661 6043 5695
rect 3188 5593 3222 5627
rect 2053 5525 2087 5559
rect 4169 5525 4203 5559
rect 3893 5321 3927 5355
rect 4813 5321 4847 5355
rect 5273 5321 5307 5355
rect 2605 5253 2639 5287
rect 1961 5185 1995 5219
rect 5181 5185 5215 5219
rect 5457 5117 5491 5151
rect 2145 4981 2179 5015
rect 2513 4777 2547 4811
rect 2973 4777 3007 4811
rect 5365 4777 5399 4811
rect 5917 4777 5951 4811
rect 1961 4709 1995 4743
rect 2053 4573 2087 4607
rect 2697 4573 2731 4607
rect 2789 4573 2823 4607
rect 3065 4573 3099 4607
rect 3985 4573 4019 4607
rect 4252 4573 4286 4607
rect 5825 4573 5859 4607
rect 5365 4233 5399 4267
rect 1869 4097 1903 4131
rect 2605 4097 2639 4131
rect 3332 4097 3366 4131
rect 5273 4097 5307 4131
rect 3065 4029 3099 4063
rect 5457 4029 5491 4063
rect 1685 3893 1719 3927
rect 2513 3893 2547 3927
rect 4445 3893 4479 3927
rect 4905 3893 4939 3927
rect 1685 3689 1719 3723
rect 2697 3689 2731 3723
rect 6561 3689 6595 3723
rect 2145 3621 2179 3655
rect 3249 3553 3283 3587
rect 4077 3553 4111 3587
rect 5181 3553 5215 3587
rect 1869 3485 1903 3519
rect 1961 3485 1995 3519
rect 2237 3485 2271 3519
rect 3157 3485 3191 3519
rect 4261 3485 4295 3519
rect 5426 3417 5460 3451
rect 3065 3349 3099 3383
rect 4353 3349 4387 3383
rect 4721 3349 4755 3383
rect 2053 3145 2087 3179
rect 4721 3145 4755 3179
rect 5365 3145 5399 3179
rect 5825 3145 5859 3179
rect 3586 3077 3620 3111
rect 2053 3009 2087 3043
rect 2605 3009 2639 3043
rect 5181 3009 5215 3043
rect 6009 3009 6043 3043
rect 2881 2941 2915 2975
rect 3341 2941 3375 2975
rect 2421 2601 2455 2635
rect 3985 2601 4019 2635
rect 4445 2601 4479 2635
rect 5181 2533 5215 2567
rect 1869 2397 1903 2431
rect 2329 2397 2363 2431
rect 3433 2397 3467 2431
rect 4169 2397 4203 2431
rect 4261 2397 4295 2431
rect 4537 2397 4571 2431
rect 4997 2397 5031 2431
rect 5733 2397 5767 2431
rect 1685 2261 1719 2295
rect 3249 2261 3283 2295
rect 5917 2261 5951 2295
<< metal1 >>
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 7282 8344 7288 8356
rect 5224 8316 7288 8344
rect 5224 8304 5230 8316
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 1104 8186 7084 8208
rect 1104 8134 1697 8186
rect 1749 8134 1761 8186
rect 1813 8134 1825 8186
rect 1877 8134 1889 8186
rect 1941 8134 1953 8186
rect 2005 8134 3192 8186
rect 3244 8134 3256 8186
rect 3308 8134 3320 8186
rect 3372 8134 3384 8186
rect 3436 8134 3448 8186
rect 3500 8134 4687 8186
rect 4739 8134 4751 8186
rect 4803 8134 4815 8186
rect 4867 8134 4879 8186
rect 4931 8134 4943 8186
rect 4995 8134 6182 8186
rect 6234 8134 6246 8186
rect 6298 8134 6310 8186
rect 6362 8134 6374 8186
rect 6426 8134 6438 8186
rect 6490 8134 7084 8186
rect 1104 8112 7084 8134
rect 5166 8032 5172 8084
rect 5224 8032 5230 8084
rect 5905 8075 5963 8081
rect 5905 8041 5917 8075
rect 5951 8072 5963 8075
rect 6086 8072 6092 8084
rect 5951 8044 6092 8072
rect 5951 8041 5963 8044
rect 5905 8035 5963 8041
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3568 7840 3985 7868
rect 3568 7828 3574 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4580 7840 4997 7868
rect 4580 7828 4586 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5224 7840 5733 7868
rect 5224 7828 5230 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 3050 7760 3056 7812
rect 3108 7800 3114 7812
rect 3329 7803 3387 7809
rect 3329 7800 3341 7803
rect 3108 7772 3341 7800
rect 3108 7760 3114 7772
rect 3329 7769 3341 7772
rect 3375 7769 3387 7803
rect 3329 7763 3387 7769
rect 2038 7692 2044 7744
rect 2096 7692 2102 7744
rect 4157 7735 4215 7741
rect 4157 7701 4169 7735
rect 4203 7732 4215 7735
rect 4430 7732 4436 7744
rect 4203 7704 4436 7732
rect 4203 7701 4215 7704
rect 4157 7695 4215 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 1104 7642 7156 7664
rect 1104 7590 2357 7642
rect 2409 7590 2421 7642
rect 2473 7590 2485 7642
rect 2537 7590 2549 7642
rect 2601 7590 2613 7642
rect 2665 7590 3852 7642
rect 3904 7590 3916 7642
rect 3968 7590 3980 7642
rect 4032 7590 4044 7642
rect 4096 7590 4108 7642
rect 4160 7590 5347 7642
rect 5399 7590 5411 7642
rect 5463 7590 5475 7642
rect 5527 7590 5539 7642
rect 5591 7590 5603 7642
rect 5655 7590 6842 7642
rect 6894 7590 6906 7642
rect 6958 7590 6970 7642
rect 7022 7590 7034 7642
rect 7086 7590 7098 7642
rect 7150 7590 7156 7642
rect 1104 7568 7156 7590
rect 934 7488 940 7540
rect 992 7528 998 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 992 7500 1685 7528
rect 992 7488 998 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 1673 7491 1731 7497
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 1872 7324 1900 7355
rect 2038 7352 2044 7404
rect 2096 7392 2102 7404
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 2096 7364 2329 7392
rect 2096 7352 2102 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2924 7364 2973 7392
rect 2924 7352 2930 7364
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 2130 7324 2136 7336
rect 1872 7296 2136 7324
rect 2130 7284 2136 7296
rect 2188 7284 2194 7336
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2096 7160 2421 7188
rect 2096 7148 2102 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2409 7151 2467 7157
rect 3050 7148 3056 7200
rect 3108 7188 3114 7200
rect 4249 7191 4307 7197
rect 4249 7188 4261 7191
rect 3108 7160 4261 7188
rect 3108 7148 3114 7160
rect 4249 7157 4261 7160
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 1104 7098 7084 7120
rect 1104 7046 1697 7098
rect 1749 7046 1761 7098
rect 1813 7046 1825 7098
rect 1877 7046 1889 7098
rect 1941 7046 1953 7098
rect 2005 7046 3192 7098
rect 3244 7046 3256 7098
rect 3308 7046 3320 7098
rect 3372 7046 3384 7098
rect 3436 7046 3448 7098
rect 3500 7046 4687 7098
rect 4739 7046 4751 7098
rect 4803 7046 4815 7098
rect 4867 7046 4879 7098
rect 4931 7046 4943 7098
rect 4995 7046 6182 7098
rect 6234 7046 6246 7098
rect 6298 7046 6310 7098
rect 6362 7046 6374 7098
rect 6426 7046 6438 7098
rect 6490 7046 7084 7098
rect 1104 7024 7084 7046
rect 2038 6808 2044 6860
rect 2096 6808 2102 6860
rect 5074 6848 5080 6860
rect 4264 6820 5080 6848
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 2866 6780 2872 6792
rect 992 6752 2872 6780
rect 992 6740 998 6752
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 4264 6789 4292 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5902 6848 5908 6860
rect 5184 6820 5908 6848
rect 5184 6792 5212 6820
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4430 6740 4436 6792
rect 4488 6740 4494 6792
rect 5166 6740 5172 6792
rect 5224 6740 5230 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 2308 6715 2366 6721
rect 2308 6681 2320 6715
rect 2354 6681 2366 6715
rect 4448 6712 4476 6740
rect 5644 6712 5672 6743
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5776 6752 5825 6780
rect 5776 6740 5782 6752
rect 5813 6749 5825 6752
rect 5859 6780 5871 6783
rect 6549 6783 6607 6789
rect 5859 6752 6408 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 4448 6684 5672 6712
rect 2308 6675 2366 6681
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2332 6644 2360 6675
rect 2280 6616 2360 6644
rect 2280 6604 2286 6616
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 3016 6616 3433 6644
rect 3016 6604 3022 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4338 6644 4344 6656
rect 4111 6616 4344 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 4982 6604 4988 6656
rect 5040 6604 5046 6656
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 6380 6653 6408 6752
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 7282 6780 7288 6792
rect 6595 6752 7288 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 5721 6647 5779 6653
rect 5721 6644 5733 6647
rect 5224 6616 5733 6644
rect 5224 6604 5230 6616
rect 5721 6613 5733 6616
rect 5767 6613 5779 6647
rect 5721 6607 5779 6613
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6613 6423 6647
rect 6365 6607 6423 6613
rect 1104 6554 7156 6576
rect 1104 6502 2357 6554
rect 2409 6502 2421 6554
rect 2473 6502 2485 6554
rect 2537 6502 2549 6554
rect 2601 6502 2613 6554
rect 2665 6502 3852 6554
rect 3904 6502 3916 6554
rect 3968 6502 3980 6554
rect 4032 6502 4044 6554
rect 4096 6502 4108 6554
rect 4160 6502 5347 6554
rect 5399 6502 5411 6554
rect 5463 6502 5475 6554
rect 5527 6502 5539 6554
rect 5591 6502 5603 6554
rect 5655 6502 6842 6554
rect 6894 6502 6906 6554
rect 6958 6502 6970 6554
rect 7022 6502 7034 6554
rect 7086 6502 7098 6554
rect 7150 6502 7156 6554
rect 1104 6480 7156 6502
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4580 6412 4629 6440
rect 4580 6400 4586 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 4982 6372 4988 6384
rect 3436 6344 4988 6372
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3436 6313 3464 6344
rect 4982 6332 4988 6344
rect 5040 6332 5046 6384
rect 3154 6307 3212 6313
rect 3154 6304 3166 6307
rect 2924 6276 3166 6304
rect 2924 6264 2930 6276
rect 3154 6273 3166 6276
rect 3200 6273 3212 6307
rect 3154 6267 3212 6273
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 3752 6276 3893 6304
rect 3752 6264 3758 6276
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 5730 6307 5788 6313
rect 5730 6304 5742 6307
rect 5316 6276 5742 6304
rect 5316 6264 5322 6276
rect 5730 6273 5742 6276
rect 5776 6273 5788 6307
rect 5730 6267 5788 6273
rect 5994 6196 6000 6248
rect 6052 6196 6058 6248
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 2130 6100 2136 6112
rect 2087 6072 2136 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3568 6072 3985 6100
rect 3568 6060 3574 6072
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 3973 6063 4031 6069
rect 1104 6010 7084 6032
rect 1104 5958 1697 6010
rect 1749 5958 1761 6010
rect 1813 5958 1825 6010
rect 1877 5958 1889 6010
rect 1941 5958 1953 6010
rect 2005 5958 3192 6010
rect 3244 5958 3256 6010
rect 3308 5958 3320 6010
rect 3372 5958 3384 6010
rect 3436 5958 3448 6010
rect 3500 5958 4687 6010
rect 4739 5958 4751 6010
rect 4803 5958 4815 6010
rect 4867 5958 4879 6010
rect 4931 5958 4943 6010
rect 4995 5958 6182 6010
rect 6234 5958 6246 6010
rect 6298 5958 6310 6010
rect 6362 5958 6374 6010
rect 6426 5958 6438 6010
rect 6490 5958 7084 6010
rect 1104 5936 7084 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 4338 5896 4344 5908
rect 1544 5868 4344 5896
rect 1544 5856 1550 5868
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5258 5856 5264 5908
rect 5316 5856 5322 5908
rect 4356 5828 4384 5856
rect 4356 5800 5028 5828
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 3510 5760 3516 5772
rect 3467 5732 3516 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4488 5732 4813 5760
rect 4488 5720 4494 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4614 5692 4620 5704
rect 4019 5664 4620 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 5000 5701 5028 5800
rect 5718 5720 5724 5772
rect 5776 5720 5782 5772
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 3176 5627 3234 5633
rect 3176 5593 3188 5627
rect 3222 5624 3234 5627
rect 3222 5596 4476 5624
rect 3222 5593 3234 5596
rect 3176 5587 3234 5593
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 1636 5528 2053 5556
rect 1636 5516 1642 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 4246 5556 4252 5568
rect 4203 5528 4252 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4448 5556 4476 5596
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 5092 5624 5120 5655
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5316 5664 6009 5692
rect 5316 5652 5322 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 4580 5596 5120 5624
rect 4580 5584 4586 5596
rect 5810 5556 5816 5568
rect 4448 5528 5816 5556
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 1104 5466 7156 5488
rect 1104 5414 2357 5466
rect 2409 5414 2421 5466
rect 2473 5414 2485 5466
rect 2537 5414 2549 5466
rect 2601 5414 2613 5466
rect 2665 5414 3852 5466
rect 3904 5414 3916 5466
rect 3968 5414 3980 5466
rect 4032 5414 4044 5466
rect 4096 5414 4108 5466
rect 4160 5414 5347 5466
rect 5399 5414 5411 5466
rect 5463 5414 5475 5466
rect 5527 5414 5539 5466
rect 5591 5414 5603 5466
rect 5655 5414 6842 5466
rect 6894 5414 6906 5466
rect 6958 5414 6970 5466
rect 7022 5414 7034 5466
rect 7086 5414 7098 5466
rect 7150 5414 7156 5466
rect 1104 5392 7156 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 3881 5355 3939 5361
rect 3881 5352 3893 5355
rect 3752 5324 3893 5352
rect 3752 5312 3758 5324
rect 3881 5321 3893 5324
rect 3927 5321 3939 5355
rect 3881 5315 3939 5321
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4672 5324 4813 5352
rect 4672 5312 4678 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 4801 5315 4859 5321
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 5224 5324 5273 5352
rect 5224 5312 5230 5324
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5284 2651 5287
rect 3050 5284 3056 5296
rect 2639 5256 3056 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2682 5216 2688 5228
rect 1995 5188 2688 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 5132 5188 5181 5216
rect 5132 5176 5138 5188
rect 5169 5185 5181 5188
rect 5215 5216 5227 5219
rect 5258 5216 5264 5228
rect 5215 5188 5264 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5408 5120 5457 5148
rect 5408 5108 5414 5120
rect 5445 5117 5457 5120
rect 5491 5148 5503 5151
rect 5902 5148 5908 5160
rect 5491 5120 5908 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 3050 5012 3056 5024
rect 2179 4984 3056 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 1104 4922 7084 4944
rect 1104 4870 1697 4922
rect 1749 4870 1761 4922
rect 1813 4870 1825 4922
rect 1877 4870 1889 4922
rect 1941 4870 1953 4922
rect 2005 4870 3192 4922
rect 3244 4870 3256 4922
rect 3308 4870 3320 4922
rect 3372 4870 3384 4922
rect 3436 4870 3448 4922
rect 3500 4870 4687 4922
rect 4739 4870 4751 4922
rect 4803 4870 4815 4922
rect 4867 4870 4879 4922
rect 4931 4870 4943 4922
rect 4995 4870 6182 4922
rect 6234 4870 6246 4922
rect 6298 4870 6310 4922
rect 6362 4870 6374 4922
rect 6426 4870 6438 4922
rect 6490 4870 7084 4922
rect 1104 4848 7084 4870
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4808 2559 4811
rect 2866 4808 2872 4820
rect 2547 4780 2872 4808
rect 2547 4777 2559 4780
rect 2501 4771 2559 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 2961 4811 3019 4817
rect 2961 4777 2973 4811
rect 3007 4808 3019 4811
rect 4614 4808 4620 4820
rect 3007 4780 4620 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4740 2007 4743
rect 2038 4740 2044 4752
rect 1995 4712 2044 4740
rect 1995 4709 2007 4712
rect 1949 4703 2007 4709
rect 2038 4700 2044 4712
rect 2096 4740 2102 4752
rect 2976 4740 3004 4771
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5350 4768 5356 4820
rect 5408 4768 5414 4820
rect 5905 4811 5963 4817
rect 5905 4777 5917 4811
rect 5951 4808 5963 4811
rect 5994 4808 6000 4820
rect 5951 4780 6000 4808
rect 5951 4777 5963 4780
rect 5905 4771 5963 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 2096 4712 3004 4740
rect 2096 4700 2102 4712
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2188 4644 2820 4672
rect 2188 4632 2194 4644
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 2792 4613 2820 4644
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 2004 4576 2053 4604
rect 2004 4564 2010 4576
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 1486 4496 1492 4548
rect 1544 4536 1550 4548
rect 2700 4536 2728 4567
rect 1544 4508 2728 4536
rect 3068 4536 3096 4567
rect 3510 4564 3516 4616
rect 3568 4604 3574 4616
rect 4246 4613 4252 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3568 4576 3985 4604
rect 3568 4564 3574 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 4240 4604 4252 4613
rect 4207 4576 4252 4604
rect 3973 4567 4031 4573
rect 4240 4567 4252 4576
rect 4246 4564 4252 4567
rect 4304 4564 4310 4616
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5132 4576 5825 4604
rect 5132 4564 5138 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5166 4536 5172 4548
rect 3068 4508 5172 4536
rect 1544 4496 1550 4508
rect 5166 4496 5172 4508
rect 5224 4496 5230 4548
rect 1104 4378 7156 4400
rect 1104 4326 2357 4378
rect 2409 4326 2421 4378
rect 2473 4326 2485 4378
rect 2537 4326 2549 4378
rect 2601 4326 2613 4378
rect 2665 4326 3852 4378
rect 3904 4326 3916 4378
rect 3968 4326 3980 4378
rect 4032 4326 4044 4378
rect 4096 4326 4108 4378
rect 4160 4326 5347 4378
rect 5399 4326 5411 4378
rect 5463 4326 5475 4378
rect 5527 4326 5539 4378
rect 5591 4326 5603 4378
rect 5655 4326 6842 4378
rect 6894 4326 6906 4378
rect 6958 4326 6970 4378
rect 7022 4326 7034 4378
rect 7086 4326 7098 4378
rect 7150 4326 7156 4378
rect 1104 4304 7156 4326
rect 1946 4224 1952 4276
rect 2004 4264 2010 4276
rect 2004 4236 2774 4264
rect 2004 4224 2010 4236
rect 2746 4196 2774 4236
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 5258 4264 5264 4276
rect 4396 4236 5264 4264
rect 4396 4224 4402 4236
rect 5258 4224 5264 4236
rect 5316 4264 5322 4276
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 5316 4236 5365 4264
rect 5316 4224 5322 4236
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 5353 4227 5411 4233
rect 2746 4168 5028 4196
rect 5000 4140 5028 4168
rect 5166 4156 5172 4208
rect 5224 4196 5230 4208
rect 5224 4168 5488 4196
rect 5224 4156 5230 4168
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2774 4128 2780 4140
rect 2639 4100 2780 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 1872 3992 1900 4091
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3320 4131 3378 4137
rect 3320 4097 3332 4131
rect 3366 4128 3378 4131
rect 3602 4128 3608 4140
rect 3366 4100 3608 4128
rect 3366 4097 3378 4100
rect 3320 4091 3378 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 5040 4100 5273 4128
rect 5040 4088 5046 4100
rect 5261 4097 5273 4100
rect 5307 4128 5319 4131
rect 5350 4128 5356 4140
rect 5307 4100 5356 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 5460 4069 5488 4168
rect 3053 4063 3111 4069
rect 3053 4060 3065 4063
rect 2096 4032 3065 4060
rect 2096 4020 2102 4032
rect 3053 4029 3065 4032
rect 3099 4029 3111 4063
rect 3053 4023 3111 4029
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5718 4060 5724 4072
rect 5491 4032 5724 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5718 4020 5724 4032
rect 5776 4060 5782 4072
rect 6546 4060 6552 4072
rect 5776 4032 6552 4060
rect 5776 4020 5782 4032
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 2958 3992 2964 4004
rect 1872 3964 2964 3992
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1673 3927 1731 3933
rect 1673 3924 1685 3927
rect 992 3896 1685 3924
rect 992 3884 998 3896
rect 1673 3893 1685 3896
rect 1719 3893 1731 3927
rect 1673 3887 1731 3893
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 4154 3924 4160 3936
rect 2547 3896 4160 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4304 3896 4445 3924
rect 4304 3884 4310 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 5166 3924 5172 3936
rect 4939 3896 5172 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 1104 3834 7084 3856
rect 1104 3782 1697 3834
rect 1749 3782 1761 3834
rect 1813 3782 1825 3834
rect 1877 3782 1889 3834
rect 1941 3782 1953 3834
rect 2005 3782 3192 3834
rect 3244 3782 3256 3834
rect 3308 3782 3320 3834
rect 3372 3782 3384 3834
rect 3436 3782 3448 3834
rect 3500 3782 4687 3834
rect 4739 3782 4751 3834
rect 4803 3782 4815 3834
rect 4867 3782 4879 3834
rect 4931 3782 4943 3834
rect 4995 3782 6182 3834
rect 6234 3782 6246 3834
rect 6298 3782 6310 3834
rect 6362 3782 6374 3834
rect 6426 3782 6438 3834
rect 6490 3782 7084 3834
rect 1104 3760 7084 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2222 3720 2228 3732
rect 1719 3692 2228 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2682 3680 2688 3732
rect 2740 3680 2746 3732
rect 5074 3720 5080 3732
rect 3252 3692 5080 3720
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 2133 3655 2191 3661
rect 2133 3652 2145 3655
rect 1636 3624 2145 3652
rect 1636 3612 1642 3624
rect 2133 3621 2145 3624
rect 2179 3652 2191 3655
rect 3252 3652 3280 3692
rect 2179 3624 3280 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 1486 3544 1492 3596
rect 1544 3584 1550 3596
rect 1544 3556 1992 3584
rect 1544 3544 1550 3556
rect 1964 3528 1992 3556
rect 2148 3528 2176 3615
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 4080 3593 4108 3692
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5350 3720 5356 3732
rect 5184 3692 5356 3720
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 5184 3652 5212 3692
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 6546 3680 6552 3732
rect 6604 3680 6610 3732
rect 4672 3624 5212 3652
rect 4672 3612 4678 3624
rect 3237 3587 3295 3593
rect 3237 3584 3249 3587
rect 2740 3556 3249 3584
rect 2740 3544 2746 3556
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 1872 3448 1900 3479
rect 1946 3476 1952 3528
rect 2004 3476 2010 3528
rect 2130 3476 2136 3528
rect 2188 3476 2194 3528
rect 2222 3476 2228 3528
rect 2280 3476 2286 3528
rect 2958 3448 2964 3460
rect 1872 3420 2964 3448
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 3068 3448 3096 3556
rect 3237 3553 3249 3556
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 4212 3556 5181 3584
rect 4212 3544 4218 3556
rect 5169 3553 5181 3556
rect 5215 3553 5227 3587
rect 5169 3547 5227 3553
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 3191 3488 4261 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 4249 3485 4261 3488
rect 4295 3516 4307 3519
rect 4338 3516 4344 3528
rect 4295 3488 4344 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4430 3448 4436 3460
rect 3068 3420 4436 3448
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5414 3451 5472 3457
rect 5414 3448 5426 3451
rect 5316 3420 5426 3448
rect 5316 3408 5322 3420
rect 5414 3417 5426 3420
rect 5460 3417 5472 3451
rect 5414 3411 5472 3417
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 4341 3383 4399 3389
rect 4341 3380 4353 3383
rect 3099 3352 4353 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 4341 3349 4353 3352
rect 4387 3380 4399 3383
rect 4614 3380 4620 3392
rect 4387 3352 4620 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4709 3383 4767 3389
rect 4709 3349 4721 3383
rect 4755 3380 4767 3383
rect 5994 3380 6000 3392
rect 4755 3352 6000 3380
rect 4755 3349 4767 3352
rect 4709 3343 4767 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 1104 3290 7156 3312
rect 1104 3238 2357 3290
rect 2409 3238 2421 3290
rect 2473 3238 2485 3290
rect 2537 3238 2549 3290
rect 2601 3238 2613 3290
rect 2665 3238 3852 3290
rect 3904 3238 3916 3290
rect 3968 3238 3980 3290
rect 4032 3238 4044 3290
rect 4096 3238 4108 3290
rect 4160 3238 5347 3290
rect 5399 3238 5411 3290
rect 5463 3238 5475 3290
rect 5527 3238 5539 3290
rect 5591 3238 5603 3290
rect 5655 3238 6842 3290
rect 6894 3238 6906 3290
rect 6958 3238 6970 3290
rect 7022 3238 7034 3290
rect 7086 3238 7098 3290
rect 7150 3238 7156 3290
rect 1104 3216 7156 3238
rect 2038 3136 2044 3188
rect 2096 3136 2102 3188
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 4488 3148 4721 3176
rect 4488 3136 4494 3148
rect 4709 3145 4721 3148
rect 4755 3145 4767 3179
rect 4709 3139 4767 3145
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 5316 3148 5365 3176
rect 5316 3136 5322 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5353 3139 5411 3145
rect 5810 3136 5816 3188
rect 5868 3136 5874 3188
rect 2314 3108 2320 3120
rect 2056 3080 2320 3108
rect 2056 3049 2084 3080
rect 2314 3068 2320 3080
rect 2372 3108 2378 3120
rect 2682 3108 2688 3120
rect 2372 3080 2688 3108
rect 2372 3068 2378 3080
rect 2682 3068 2688 3080
rect 2740 3068 2746 3120
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 3574 3111 3632 3117
rect 3574 3108 3586 3111
rect 3108 3080 3586 3108
rect 3108 3068 3114 3080
rect 3574 3077 3586 3080
rect 3620 3077 3632 3111
rect 3574 3071 3632 3077
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2188 3012 2605 3040
rect 2188 3000 2194 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 5166 3000 5172 3052
rect 5224 3000 5230 3052
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 2915 2944 3341 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 4246 2836 4252 2848
rect 2004 2808 4252 2836
rect 2004 2796 2010 2808
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 1104 2746 7084 2768
rect 1104 2694 1697 2746
rect 1749 2694 1761 2746
rect 1813 2694 1825 2746
rect 1877 2694 1889 2746
rect 1941 2694 1953 2746
rect 2005 2694 3192 2746
rect 3244 2694 3256 2746
rect 3308 2694 3320 2746
rect 3372 2694 3384 2746
rect 3436 2694 3448 2746
rect 3500 2694 4687 2746
rect 4739 2694 4751 2746
rect 4803 2694 4815 2746
rect 4867 2694 4879 2746
rect 4931 2694 4943 2746
rect 4995 2694 6182 2746
rect 6234 2694 6246 2746
rect 6298 2694 6310 2746
rect 6362 2694 6374 2746
rect 6426 2694 6438 2746
rect 6490 2694 7084 2746
rect 1104 2672 7084 2694
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 3510 2632 3516 2644
rect 2455 2604 3516 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3660 2604 3985 2632
rect 3660 2592 3666 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 5902 2632 5908 2644
rect 4479 2604 5908 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 4448 2564 4476 2595
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 2832 2536 4476 2564
rect 5169 2567 5227 2573
rect 2832 2524 2838 2536
rect 5169 2533 5181 2567
rect 5215 2564 5227 2567
rect 7282 2564 7288 2576
rect 5215 2536 7288 2564
rect 5215 2533 5227 2536
rect 5169 2527 5227 2533
rect 7282 2524 7288 2536
rect 7340 2524 7346 2576
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2314 2428 2320 2440
rect 1903 2400 2320 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4154 2428 4160 2440
rect 3467 2400 4160 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4246 2388 4252 2440
rect 4304 2388 4310 2440
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5074 2428 5080 2440
rect 5031 2400 5080 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5074 2388 5080 2400
rect 5132 2388 5138 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 72 2264 1685 2292
rect 72 2252 78 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2252 3298 2304
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 6454 2292 6460 2304
rect 5951 2264 6460 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 1104 2202 7156 2224
rect 1104 2150 2357 2202
rect 2409 2150 2421 2202
rect 2473 2150 2485 2202
rect 2537 2150 2549 2202
rect 2601 2150 2613 2202
rect 2665 2150 3852 2202
rect 3904 2150 3916 2202
rect 3968 2150 3980 2202
rect 4032 2150 4044 2202
rect 4096 2150 4108 2202
rect 4160 2150 5347 2202
rect 5399 2150 5411 2202
rect 5463 2150 5475 2202
rect 5527 2150 5539 2202
rect 5591 2150 5603 2202
rect 5655 2150 6842 2202
rect 6894 2150 6906 2202
rect 6958 2150 6970 2202
rect 7022 2150 7034 2202
rect 7086 2150 7098 2202
rect 7150 2150 7156 2202
rect 1104 2128 7156 2150
<< via1 >>
rect 5172 8304 5224 8356
rect 7288 8304 7340 8356
rect 1697 8134 1749 8186
rect 1761 8134 1813 8186
rect 1825 8134 1877 8186
rect 1889 8134 1941 8186
rect 1953 8134 2005 8186
rect 3192 8134 3244 8186
rect 3256 8134 3308 8186
rect 3320 8134 3372 8186
rect 3384 8134 3436 8186
rect 3448 8134 3500 8186
rect 4687 8134 4739 8186
rect 4751 8134 4803 8186
rect 4815 8134 4867 8186
rect 4879 8134 4931 8186
rect 4943 8134 4995 8186
rect 6182 8134 6234 8186
rect 6246 8134 6298 8186
rect 6310 8134 6362 8186
rect 6374 8134 6426 8186
rect 6438 8134 6490 8186
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 6092 8032 6144 8084
rect 3516 7828 3568 7880
rect 4528 7828 4580 7880
rect 5172 7828 5224 7880
rect 3056 7760 3108 7812
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 4436 7692 4488 7744
rect 2357 7590 2409 7642
rect 2421 7590 2473 7642
rect 2485 7590 2537 7642
rect 2549 7590 2601 7642
rect 2613 7590 2665 7642
rect 3852 7590 3904 7642
rect 3916 7590 3968 7642
rect 3980 7590 4032 7642
rect 4044 7590 4096 7642
rect 4108 7590 4160 7642
rect 5347 7590 5399 7642
rect 5411 7590 5463 7642
rect 5475 7590 5527 7642
rect 5539 7590 5591 7642
rect 5603 7590 5655 7642
rect 6842 7590 6894 7642
rect 6906 7590 6958 7642
rect 6970 7590 7022 7642
rect 7034 7590 7086 7642
rect 7098 7590 7150 7642
rect 940 7488 992 7540
rect 2044 7352 2096 7404
rect 2872 7352 2924 7404
rect 2136 7284 2188 7336
rect 2044 7148 2096 7200
rect 3056 7148 3108 7200
rect 1697 7046 1749 7098
rect 1761 7046 1813 7098
rect 1825 7046 1877 7098
rect 1889 7046 1941 7098
rect 1953 7046 2005 7098
rect 3192 7046 3244 7098
rect 3256 7046 3308 7098
rect 3320 7046 3372 7098
rect 3384 7046 3436 7098
rect 3448 7046 3500 7098
rect 4687 7046 4739 7098
rect 4751 7046 4803 7098
rect 4815 7046 4867 7098
rect 4879 7046 4931 7098
rect 4943 7046 4995 7098
rect 6182 7046 6234 7098
rect 6246 7046 6298 7098
rect 6310 7046 6362 7098
rect 6374 7046 6426 7098
rect 6438 7046 6490 7098
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 940 6740 992 6792
rect 2872 6740 2924 6792
rect 5080 6808 5132 6860
rect 5908 6808 5960 6860
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5724 6740 5776 6792
rect 2228 6604 2280 6656
rect 2964 6604 3016 6656
rect 4344 6604 4396 6656
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 5172 6604 5224 6656
rect 7288 6740 7340 6792
rect 2357 6502 2409 6554
rect 2421 6502 2473 6554
rect 2485 6502 2537 6554
rect 2549 6502 2601 6554
rect 2613 6502 2665 6554
rect 3852 6502 3904 6554
rect 3916 6502 3968 6554
rect 3980 6502 4032 6554
rect 4044 6502 4096 6554
rect 4108 6502 4160 6554
rect 5347 6502 5399 6554
rect 5411 6502 5463 6554
rect 5475 6502 5527 6554
rect 5539 6502 5591 6554
rect 5603 6502 5655 6554
rect 6842 6502 6894 6554
rect 6906 6502 6958 6554
rect 6970 6502 7022 6554
rect 7034 6502 7086 6554
rect 7098 6502 7150 6554
rect 4528 6400 4580 6452
rect 2872 6264 2924 6316
rect 4988 6332 5040 6384
rect 3700 6264 3752 6316
rect 5264 6264 5316 6316
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 2136 6060 2188 6112
rect 3516 6060 3568 6112
rect 1697 5958 1749 6010
rect 1761 5958 1813 6010
rect 1825 5958 1877 6010
rect 1889 5958 1941 6010
rect 1953 5958 2005 6010
rect 3192 5958 3244 6010
rect 3256 5958 3308 6010
rect 3320 5958 3372 6010
rect 3384 5958 3436 6010
rect 3448 5958 3500 6010
rect 4687 5958 4739 6010
rect 4751 5958 4803 6010
rect 4815 5958 4867 6010
rect 4879 5958 4931 6010
rect 4943 5958 4995 6010
rect 6182 5958 6234 6010
rect 6246 5958 6298 6010
rect 6310 5958 6362 6010
rect 6374 5958 6426 6010
rect 6438 5958 6490 6010
rect 1492 5856 1544 5908
rect 4344 5856 4396 5908
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 3516 5720 3568 5772
rect 4436 5720 4488 5772
rect 4620 5652 4672 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 5724 5763 5776 5772
rect 5724 5729 5733 5763
rect 5733 5729 5767 5763
rect 5767 5729 5776 5763
rect 5724 5720 5776 5729
rect 1584 5516 1636 5568
rect 4252 5516 4304 5568
rect 4528 5584 4580 5636
rect 5264 5652 5316 5704
rect 5816 5516 5868 5568
rect 2357 5414 2409 5466
rect 2421 5414 2473 5466
rect 2485 5414 2537 5466
rect 2549 5414 2601 5466
rect 2613 5414 2665 5466
rect 3852 5414 3904 5466
rect 3916 5414 3968 5466
rect 3980 5414 4032 5466
rect 4044 5414 4096 5466
rect 4108 5414 4160 5466
rect 5347 5414 5399 5466
rect 5411 5414 5463 5466
rect 5475 5414 5527 5466
rect 5539 5414 5591 5466
rect 5603 5414 5655 5466
rect 6842 5414 6894 5466
rect 6906 5414 6958 5466
rect 6970 5414 7022 5466
rect 7034 5414 7086 5466
rect 7098 5414 7150 5466
rect 3700 5312 3752 5364
rect 4620 5312 4672 5364
rect 5172 5312 5224 5364
rect 3056 5244 3108 5296
rect 2688 5176 2740 5228
rect 5080 5176 5132 5228
rect 5264 5176 5316 5228
rect 5356 5108 5408 5160
rect 5908 5108 5960 5160
rect 3056 4972 3108 5024
rect 1697 4870 1749 4922
rect 1761 4870 1813 4922
rect 1825 4870 1877 4922
rect 1889 4870 1941 4922
rect 1953 4870 2005 4922
rect 3192 4870 3244 4922
rect 3256 4870 3308 4922
rect 3320 4870 3372 4922
rect 3384 4870 3436 4922
rect 3448 4870 3500 4922
rect 4687 4870 4739 4922
rect 4751 4870 4803 4922
rect 4815 4870 4867 4922
rect 4879 4870 4931 4922
rect 4943 4870 4995 4922
rect 6182 4870 6234 4922
rect 6246 4870 6298 4922
rect 6310 4870 6362 4922
rect 6374 4870 6426 4922
rect 6438 4870 6490 4922
rect 2872 4768 2924 4820
rect 2044 4700 2096 4752
rect 4620 4768 4672 4820
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 6000 4768 6052 4820
rect 2136 4632 2188 4684
rect 1952 4564 2004 4616
rect 1492 4496 1544 4548
rect 3516 4564 3568 4616
rect 4252 4607 4304 4616
rect 4252 4573 4286 4607
rect 4286 4573 4304 4607
rect 4252 4564 4304 4573
rect 5080 4564 5132 4616
rect 5172 4496 5224 4548
rect 2357 4326 2409 4378
rect 2421 4326 2473 4378
rect 2485 4326 2537 4378
rect 2549 4326 2601 4378
rect 2613 4326 2665 4378
rect 3852 4326 3904 4378
rect 3916 4326 3968 4378
rect 3980 4326 4032 4378
rect 4044 4326 4096 4378
rect 4108 4326 4160 4378
rect 5347 4326 5399 4378
rect 5411 4326 5463 4378
rect 5475 4326 5527 4378
rect 5539 4326 5591 4378
rect 5603 4326 5655 4378
rect 6842 4326 6894 4378
rect 6906 4326 6958 4378
rect 6970 4326 7022 4378
rect 7034 4326 7086 4378
rect 7098 4326 7150 4378
rect 1952 4224 2004 4276
rect 4344 4224 4396 4276
rect 5264 4224 5316 4276
rect 5172 4156 5224 4208
rect 2780 4088 2832 4140
rect 3608 4088 3660 4140
rect 4988 4088 5040 4140
rect 5356 4088 5408 4140
rect 2044 4020 2096 4072
rect 5724 4020 5776 4072
rect 6552 4020 6604 4072
rect 2964 3952 3016 4004
rect 940 3884 992 3936
rect 4160 3884 4212 3936
rect 4252 3884 4304 3936
rect 5172 3884 5224 3936
rect 1697 3782 1749 3834
rect 1761 3782 1813 3834
rect 1825 3782 1877 3834
rect 1889 3782 1941 3834
rect 1953 3782 2005 3834
rect 3192 3782 3244 3834
rect 3256 3782 3308 3834
rect 3320 3782 3372 3834
rect 3384 3782 3436 3834
rect 3448 3782 3500 3834
rect 4687 3782 4739 3834
rect 4751 3782 4803 3834
rect 4815 3782 4867 3834
rect 4879 3782 4931 3834
rect 4943 3782 4995 3834
rect 6182 3782 6234 3834
rect 6246 3782 6298 3834
rect 6310 3782 6362 3834
rect 6374 3782 6426 3834
rect 6438 3782 6490 3834
rect 2228 3680 2280 3732
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 1584 3612 1636 3664
rect 1492 3544 1544 3596
rect 2688 3544 2740 3596
rect 5080 3680 5132 3732
rect 4620 3612 4672 3664
rect 5356 3680 5408 3732
rect 6552 3723 6604 3732
rect 6552 3689 6561 3723
rect 6561 3689 6595 3723
rect 6595 3689 6604 3723
rect 6552 3680 6604 3689
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 2136 3476 2188 3528
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 2964 3408 3016 3460
rect 4160 3544 4212 3596
rect 4344 3476 4396 3528
rect 4436 3408 4488 3460
rect 5264 3408 5316 3460
rect 4620 3340 4672 3392
rect 6000 3340 6052 3392
rect 2357 3238 2409 3290
rect 2421 3238 2473 3290
rect 2485 3238 2537 3290
rect 2549 3238 2601 3290
rect 2613 3238 2665 3290
rect 3852 3238 3904 3290
rect 3916 3238 3968 3290
rect 3980 3238 4032 3290
rect 4044 3238 4096 3290
rect 4108 3238 4160 3290
rect 5347 3238 5399 3290
rect 5411 3238 5463 3290
rect 5475 3238 5527 3290
rect 5539 3238 5591 3290
rect 5603 3238 5655 3290
rect 6842 3238 6894 3290
rect 6906 3238 6958 3290
rect 6970 3238 7022 3290
rect 7034 3238 7086 3290
rect 7098 3238 7150 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 4436 3136 4488 3188
rect 5264 3136 5316 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 2320 3068 2372 3120
rect 2688 3068 2740 3120
rect 3056 3068 3108 3120
rect 2136 3000 2188 3052
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 1952 2796 2004 2848
rect 4252 2796 4304 2848
rect 1697 2694 1749 2746
rect 1761 2694 1813 2746
rect 1825 2694 1877 2746
rect 1889 2694 1941 2746
rect 1953 2694 2005 2746
rect 3192 2694 3244 2746
rect 3256 2694 3308 2746
rect 3320 2694 3372 2746
rect 3384 2694 3436 2746
rect 3448 2694 3500 2746
rect 4687 2694 4739 2746
rect 4751 2694 4803 2746
rect 4815 2694 4867 2746
rect 4879 2694 4931 2746
rect 4943 2694 4995 2746
rect 6182 2694 6234 2746
rect 6246 2694 6298 2746
rect 6310 2694 6362 2746
rect 6374 2694 6426 2746
rect 6438 2694 6490 2746
rect 3516 2592 3568 2644
rect 3608 2592 3660 2644
rect 2780 2524 2832 2576
rect 5908 2592 5960 2644
rect 7288 2524 7340 2576
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 5080 2388 5132 2440
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 20 2252 72 2304
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 6460 2252 6512 2304
rect 2357 2150 2409 2202
rect 2421 2150 2473 2202
rect 2485 2150 2537 2202
rect 2549 2150 2601 2202
rect 2613 2150 2665 2202
rect 3852 2150 3904 2202
rect 3916 2150 3968 2202
rect 3980 2150 4032 2202
rect 4044 2150 4096 2202
rect 4108 2150 4160 2202
rect 5347 2150 5399 2202
rect 5411 2150 5463 2202
rect 5475 2150 5527 2202
rect 5539 2150 5591 2202
rect 5603 2150 5655 2202
rect 6842 2150 6894 2202
rect 6906 2150 6958 2202
rect 6970 2150 7022 2202
rect 7034 2150 7086 2202
rect 7098 2150 7150 2202
<< metal2 >>
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 952 7546 980 10231
rect 3238 9738 3294 10402
rect 6458 9738 6514 10402
rect 3238 9710 3556 9738
rect 3238 9602 3294 9710
rect 1697 8188 2005 8197
rect 1697 8186 1703 8188
rect 1759 8186 1783 8188
rect 1839 8186 1863 8188
rect 1919 8186 1943 8188
rect 1999 8186 2005 8188
rect 1759 8134 1761 8186
rect 1941 8134 1943 8186
rect 1697 8132 1703 8134
rect 1759 8132 1783 8134
rect 1839 8132 1863 8134
rect 1919 8132 1943 8134
rect 1999 8132 2005 8134
rect 1697 8123 2005 8132
rect 3192 8188 3500 8197
rect 3192 8186 3198 8188
rect 3254 8186 3278 8188
rect 3334 8186 3358 8188
rect 3414 8186 3438 8188
rect 3494 8186 3500 8188
rect 3254 8134 3256 8186
rect 3436 8134 3438 8186
rect 3192 8132 3198 8134
rect 3254 8132 3278 8134
rect 3334 8132 3358 8134
rect 3414 8132 3438 8134
rect 3494 8132 3500 8134
rect 3192 8123 3500 8132
rect 3528 7886 3556 9710
rect 6104 9710 6514 9738
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 4687 8188 4995 8197
rect 4687 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4933 8188
rect 4989 8186 4995 8188
rect 4749 8134 4751 8186
rect 4931 8134 4933 8186
rect 4687 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4933 8134
rect 4989 8132 4995 8134
rect 4687 8123 4995 8132
rect 5184 8090 5212 8298
rect 6104 8090 6132 9710
rect 6458 9602 6514 9710
rect 7286 8936 7342 8945
rect 7286 8871 7342 8880
rect 7300 8362 7328 8871
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 6182 8188 6490 8197
rect 6182 8186 6188 8188
rect 6244 8186 6268 8188
rect 6324 8186 6348 8188
rect 6404 8186 6428 8188
rect 6484 8186 6490 8188
rect 6244 8134 6246 8186
rect 6426 8134 6428 8186
rect 6182 8132 6188 8134
rect 6244 8132 6268 8134
rect 6324 8132 6348 8134
rect 6404 8132 6428 8134
rect 6484 8132 6490 8134
rect 6182 8123 6490 8132
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 940 7540 992 7546
rect 940 7482 992 7488
rect 2056 7410 2084 7686
rect 2357 7644 2665 7653
rect 2357 7642 2363 7644
rect 2419 7642 2443 7644
rect 2499 7642 2523 7644
rect 2579 7642 2603 7644
rect 2659 7642 2665 7644
rect 2419 7590 2421 7642
rect 2601 7590 2603 7642
rect 2357 7588 2363 7590
rect 2419 7588 2443 7590
rect 2499 7588 2523 7590
rect 2579 7588 2603 7590
rect 2659 7588 2665 7590
rect 2357 7579 2665 7588
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1697 7100 2005 7109
rect 1697 7098 1703 7100
rect 1759 7098 1783 7100
rect 1839 7098 1863 7100
rect 1919 7098 1943 7100
rect 1999 7098 2005 7100
rect 1759 7046 1761 7098
rect 1941 7046 1943 7098
rect 1697 7044 1703 7046
rect 1759 7044 1783 7046
rect 1839 7044 1863 7046
rect 1919 7044 1943 7046
rect 1999 7044 2005 7046
rect 1697 7035 2005 7044
rect 938 6896 994 6905
rect 2056 6866 2084 7142
rect 938 6831 994 6840
rect 2044 6860 2096 6866
rect 952 6798 980 6831
rect 2044 6802 2096 6808
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 2148 6118 2176 7278
rect 2884 6798 2912 7346
rect 3068 7206 3096 7754
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 3852 7644 4160 7653
rect 3852 7642 3858 7644
rect 3914 7642 3938 7644
rect 3994 7642 4018 7644
rect 4074 7642 4098 7644
rect 4154 7642 4160 7644
rect 3914 7590 3916 7642
rect 4096 7590 4098 7642
rect 3852 7588 3858 7590
rect 3914 7588 3938 7590
rect 3994 7588 4018 7590
rect 4074 7588 4098 7590
rect 4154 7588 4160 7590
rect 3852 7579 4160 7588
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 1697 6012 2005 6021
rect 1697 6010 1703 6012
rect 1759 6010 1783 6012
rect 1839 6010 1863 6012
rect 1919 6010 1943 6012
rect 1999 6010 2005 6012
rect 1759 5958 1761 6010
rect 1941 5958 1943 6010
rect 1697 5956 1703 5958
rect 1759 5956 1783 5958
rect 1839 5956 1863 5958
rect 1919 5956 1943 5958
rect 1999 5956 2005 5958
rect 1697 5947 2005 5956
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1504 4554 1532 5850
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 952 3505 980 3878
rect 1504 3602 1532 4490
rect 1596 3670 1624 5510
rect 1697 4924 2005 4933
rect 1697 4922 1703 4924
rect 1759 4922 1783 4924
rect 1839 4922 1863 4924
rect 1919 4922 1943 4924
rect 1999 4922 2005 4924
rect 1759 4870 1761 4922
rect 1941 4870 1943 4922
rect 1697 4868 1703 4870
rect 1759 4868 1783 4870
rect 1839 4868 1863 4870
rect 1919 4868 1943 4870
rect 1999 4868 2005 4870
rect 1697 4859 2005 4868
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 4282 1992 4558
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 2056 4162 2084 4694
rect 2148 4690 2176 6054
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2056 4134 2176 4162
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 1697 3836 2005 3845
rect 1697 3834 1703 3836
rect 1759 3834 1783 3836
rect 1839 3834 1863 3836
rect 1919 3834 1943 3836
rect 1999 3834 2005 3836
rect 1759 3782 1761 3834
rect 1941 3782 1943 3834
rect 1697 3780 1703 3782
rect 1759 3780 1783 3782
rect 1839 3780 1863 3782
rect 1919 3780 1943 3782
rect 1999 3780 2005 3782
rect 1697 3771 2005 3780
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1952 3528 2004 3534
rect 938 3496 994 3505
rect 1952 3470 2004 3476
rect 938 3431 994 3440
rect 1964 2854 1992 3470
rect 2056 3194 2084 4014
rect 2148 3618 2176 4134
rect 2240 3738 2268 6598
rect 2357 6556 2665 6565
rect 2357 6554 2363 6556
rect 2419 6554 2443 6556
rect 2499 6554 2523 6556
rect 2579 6554 2603 6556
rect 2659 6554 2665 6556
rect 2419 6502 2421 6554
rect 2601 6502 2603 6554
rect 2357 6500 2363 6502
rect 2419 6500 2443 6502
rect 2499 6500 2523 6502
rect 2579 6500 2603 6502
rect 2659 6500 2665 6502
rect 2357 6491 2665 6500
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2357 5468 2665 5477
rect 2357 5466 2363 5468
rect 2419 5466 2443 5468
rect 2499 5466 2523 5468
rect 2579 5466 2603 5468
rect 2659 5466 2665 5468
rect 2419 5414 2421 5466
rect 2601 5414 2603 5466
rect 2357 5412 2363 5414
rect 2419 5412 2443 5414
rect 2499 5412 2523 5414
rect 2579 5412 2603 5414
rect 2659 5412 2665 5414
rect 2357 5403 2665 5412
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2357 4380 2665 4389
rect 2357 4378 2363 4380
rect 2419 4378 2443 4380
rect 2499 4378 2523 4380
rect 2579 4378 2603 4380
rect 2659 4378 2665 4380
rect 2419 4326 2421 4378
rect 2601 4326 2603 4378
rect 2357 4324 2363 4326
rect 2419 4324 2443 4326
rect 2499 4324 2523 4326
rect 2579 4324 2603 4326
rect 2659 4324 2665 4326
rect 2357 4315 2665 4324
rect 2700 3738 2728 5170
rect 2884 4826 2912 6258
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2148 3590 2268 3618
rect 2240 3534 2268 3590
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2148 3058 2176 3470
rect 2357 3292 2665 3301
rect 2357 3290 2363 3292
rect 2419 3290 2443 3292
rect 2499 3290 2523 3292
rect 2579 3290 2603 3292
rect 2659 3290 2665 3292
rect 2419 3238 2421 3290
rect 2601 3238 2603 3290
rect 2357 3236 2363 3238
rect 2419 3236 2443 3238
rect 2499 3236 2523 3238
rect 2579 3236 2603 3238
rect 2659 3236 2665 3238
rect 2357 3227 2665 3236
rect 2700 3126 2728 3538
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1697 2748 2005 2757
rect 1697 2746 1703 2748
rect 1759 2746 1783 2748
rect 1839 2746 1863 2748
rect 1919 2746 1943 2748
rect 1999 2746 2005 2748
rect 1759 2694 1761 2746
rect 1941 2694 1943 2746
rect 1697 2692 1703 2694
rect 1759 2692 1783 2694
rect 1839 2692 1863 2694
rect 1919 2692 1943 2694
rect 1999 2692 2005 2694
rect 1697 2683 2005 2692
rect 2332 2446 2360 3062
rect 2792 2582 2820 4082
rect 2976 4010 3004 6598
rect 3068 5302 3096 7142
rect 3192 7100 3500 7109
rect 3192 7098 3198 7100
rect 3254 7098 3278 7100
rect 3334 7098 3358 7100
rect 3414 7098 3438 7100
rect 3494 7098 3500 7100
rect 3254 7046 3256 7098
rect 3436 7046 3438 7098
rect 3192 7044 3198 7046
rect 3254 7044 3278 7046
rect 3334 7044 3358 7046
rect 3414 7044 3438 7046
rect 3494 7044 3500 7046
rect 3192 7035 3500 7044
rect 4448 6798 4476 7686
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 3852 6556 4160 6565
rect 3852 6554 3858 6556
rect 3914 6554 3938 6556
rect 3994 6554 4018 6556
rect 4074 6554 4098 6556
rect 4154 6554 4160 6556
rect 3914 6502 3916 6554
rect 4096 6502 4098 6554
rect 3852 6500 3858 6502
rect 3914 6500 3938 6502
rect 3994 6500 4018 6502
rect 4074 6500 4098 6502
rect 4154 6500 4160 6502
rect 3852 6491 4160 6500
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3192 6012 3500 6021
rect 3192 6010 3198 6012
rect 3254 6010 3278 6012
rect 3334 6010 3358 6012
rect 3414 6010 3438 6012
rect 3494 6010 3500 6012
rect 3254 5958 3256 6010
rect 3436 5958 3438 6010
rect 3192 5956 3198 5958
rect 3254 5956 3278 5958
rect 3334 5956 3358 5958
rect 3414 5956 3438 5958
rect 3494 5956 3500 5958
rect 3192 5947 3500 5956
rect 3528 5778 3556 6054
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3712 5370 3740 6258
rect 4356 5914 4384 6598
rect 4540 6458 4568 7822
rect 4687 7100 4995 7109
rect 4687 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4933 7100
rect 4989 7098 4995 7100
rect 4749 7046 4751 7098
rect 4931 7046 4933 7098
rect 4687 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4933 7046
rect 4989 7044 4995 7046
rect 4687 7035 4995 7044
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3852 5468 4160 5477
rect 3852 5466 3858 5468
rect 3914 5466 3938 5468
rect 3994 5466 4018 5468
rect 4074 5466 4098 5468
rect 4154 5466 4160 5468
rect 3914 5414 3916 5466
rect 4096 5414 4098 5466
rect 3852 5412 3858 5414
rect 3914 5412 3938 5414
rect 3994 5412 4018 5414
rect 4074 5412 4098 5414
rect 4154 5412 4160 5414
rect 3852 5403 4160 5412
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2976 3466 3004 3946
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 3068 3126 3096 4966
rect 3192 4924 3500 4933
rect 3192 4922 3198 4924
rect 3254 4922 3278 4924
rect 3334 4922 3358 4924
rect 3414 4922 3438 4924
rect 3494 4922 3500 4924
rect 3254 4870 3256 4922
rect 3436 4870 3438 4922
rect 3192 4868 3198 4870
rect 3254 4868 3278 4870
rect 3334 4868 3358 4870
rect 3414 4868 3438 4870
rect 3494 4868 3500 4870
rect 3192 4859 3500 4868
rect 4264 4622 4292 5510
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3192 3836 3500 3845
rect 3192 3834 3198 3836
rect 3254 3834 3278 3836
rect 3334 3834 3358 3836
rect 3414 3834 3438 3836
rect 3494 3834 3500 3836
rect 3254 3782 3256 3834
rect 3436 3782 3438 3834
rect 3192 3780 3198 3782
rect 3254 3780 3278 3782
rect 3334 3780 3358 3782
rect 3414 3780 3438 3782
rect 3494 3780 3500 3782
rect 3192 3771 3500 3780
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3192 2748 3500 2757
rect 3192 2746 3198 2748
rect 3254 2746 3278 2748
rect 3334 2746 3358 2748
rect 3414 2746 3438 2748
rect 3494 2746 3500 2748
rect 3254 2694 3256 2746
rect 3436 2694 3438 2746
rect 3192 2692 3198 2694
rect 3254 2692 3278 2694
rect 3334 2692 3358 2694
rect 3414 2692 3438 2694
rect 3494 2692 3500 2694
rect 3192 2683 3500 2692
rect 3528 2650 3556 4558
rect 3852 4380 4160 4389
rect 3852 4378 3858 4380
rect 3914 4378 3938 4380
rect 3994 4378 4018 4380
rect 4074 4378 4098 4380
rect 4154 4378 4160 4380
rect 3914 4326 3916 4378
rect 4096 4326 4098 4378
rect 3852 4324 3858 4326
rect 3914 4324 3938 4326
rect 3994 4324 4018 4326
rect 4074 4324 4098 4326
rect 4154 4324 4160 4326
rect 3852 4315 4160 4324
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 2650 3648 4082
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4172 3602 4200 3878
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3852 3292 4160 3301
rect 3852 3290 3858 3292
rect 3914 3290 3938 3292
rect 3994 3290 4018 3292
rect 4074 3290 4098 3292
rect 4154 3290 4160 3292
rect 3914 3238 3916 3290
rect 4096 3238 4098 3290
rect 3852 3236 3858 3238
rect 3914 3236 3938 3238
rect 3994 3236 4018 3238
rect 4074 3236 4098 3238
rect 4154 3236 4160 3238
rect 3852 3227 4160 3236
rect 4264 3108 4292 3878
rect 4356 3534 4384 4218
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4448 3466 4476 5714
rect 4540 5642 4568 6394
rect 5000 6390 5028 6598
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4687 6012 4995 6021
rect 4687 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4933 6012
rect 4989 6010 4995 6012
rect 4749 5958 4751 6010
rect 4931 5958 4933 6010
rect 4687 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4933 5958
rect 4989 5956 4995 5958
rect 4687 5947 4995 5956
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4632 5370 4660 5646
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4724 5114 4752 5646
rect 5092 5234 5120 6802
rect 5184 6798 5212 7822
rect 5347 7644 5655 7653
rect 5347 7642 5353 7644
rect 5409 7642 5433 7644
rect 5489 7642 5513 7644
rect 5569 7642 5593 7644
rect 5649 7642 5655 7644
rect 5409 7590 5411 7642
rect 5591 7590 5593 7642
rect 5347 7588 5353 7590
rect 5409 7588 5433 7590
rect 5489 7588 5513 7590
rect 5569 7588 5593 7590
rect 5649 7588 5655 7590
rect 5347 7579 5655 7588
rect 6842 7644 7150 7653
rect 6842 7642 6848 7644
rect 6904 7642 6928 7644
rect 6984 7642 7008 7644
rect 7064 7642 7088 7644
rect 7144 7642 7150 7644
rect 6904 7590 6906 7642
rect 7086 7590 7088 7642
rect 6842 7588 6848 7590
rect 6904 7588 6928 7590
rect 6984 7588 7008 7590
rect 7064 7588 7088 7590
rect 7144 7588 7150 7590
rect 6842 7579 7150 7588
rect 6182 7100 6490 7109
rect 6182 7098 6188 7100
rect 6244 7098 6268 7100
rect 6324 7098 6348 7100
rect 6404 7098 6428 7100
rect 6484 7098 6490 7100
rect 6244 7046 6246 7098
rect 6426 7046 6428 7098
rect 6182 7044 6188 7046
rect 6244 7044 6268 7046
rect 6324 7044 6348 7046
rect 6404 7044 6428 7046
rect 6484 7044 6490 7046
rect 6182 7035 6490 7044
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 5370 5212 6598
rect 5347 6556 5655 6565
rect 5347 6554 5353 6556
rect 5409 6554 5433 6556
rect 5489 6554 5513 6556
rect 5569 6554 5593 6556
rect 5649 6554 5655 6556
rect 5409 6502 5411 6554
rect 5591 6502 5593 6554
rect 5347 6500 5353 6502
rect 5409 6500 5433 6502
rect 5489 6500 5513 6502
rect 5569 6500 5593 6502
rect 5649 6500 5655 6502
rect 5347 6491 5655 6500
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5914 5304 6258
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5736 5778 5764 6734
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4540 5086 4752 5114
rect 4540 4842 4568 5086
rect 4687 4924 4995 4933
rect 4687 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4933 4924
rect 4989 4922 4995 4924
rect 4749 4870 4751 4922
rect 4931 4870 4933 4922
rect 4687 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4933 4870
rect 4989 4868 4995 4870
rect 4687 4859 4995 4868
rect 4540 4826 4660 4842
rect 4540 4820 4672 4826
rect 4540 4814 4620 4820
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4448 3194 4476 3402
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4172 3080 4292 3108
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 4172 2446 4200 3080
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2446 4292 2790
rect 4540 2446 4568 4814
rect 4620 4762 4672 4768
rect 5092 4706 5120 5170
rect 5000 4678 5120 4706
rect 5184 4706 5212 5306
rect 5276 5234 5304 5646
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5347 5468 5655 5477
rect 5347 5466 5353 5468
rect 5409 5466 5433 5468
rect 5489 5466 5513 5468
rect 5569 5466 5593 5468
rect 5649 5466 5655 5468
rect 5409 5414 5411 5466
rect 5591 5414 5593 5466
rect 5347 5412 5353 5414
rect 5409 5412 5433 5414
rect 5489 5412 5513 5414
rect 5569 5412 5593 5414
rect 5649 5412 5655 5414
rect 5347 5403 5655 5412
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4826 5396 5102
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5184 4678 5304 4706
rect 5000 4146 5028 4678
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4687 3836 4995 3845
rect 4687 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4933 3836
rect 4989 3834 4995 3836
rect 4749 3782 4751 3834
rect 4931 3782 4933 3834
rect 4687 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4933 3782
rect 4989 3780 4995 3782
rect 4687 3771 4995 3780
rect 5092 3738 5120 4558
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5184 4214 5212 4490
rect 5276 4282 5304 4678
rect 5347 4380 5655 4389
rect 5347 4378 5353 4380
rect 5409 4378 5433 4380
rect 5489 4378 5513 4380
rect 5569 4378 5593 4380
rect 5649 4378 5655 4380
rect 5409 4326 5411 4378
rect 5591 4326 5593 4378
rect 5347 4324 5353 4326
rect 5409 4324 5433 4326
rect 5489 4324 5513 4326
rect 5569 4324 5593 4326
rect 5649 4324 5655 4326
rect 5347 4315 5655 4324
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4632 3398 4660 3606
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4687 2748 4995 2757
rect 4687 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4933 2748
rect 4989 2746 4995 2748
rect 4749 2694 4751 2746
rect 4931 2694 4933 2746
rect 4687 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4933 2694
rect 4989 2692 4995 2694
rect 4687 2683 4995 2692
rect 5092 2446 5120 3674
rect 5184 3058 5212 3878
rect 5368 3738 5396 4082
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 3194 5304 3402
rect 5347 3292 5655 3301
rect 5347 3290 5353 3292
rect 5409 3290 5433 3292
rect 5489 3290 5513 3292
rect 5569 3290 5593 3292
rect 5649 3290 5655 3292
rect 5409 3238 5411 3290
rect 5591 3238 5593 3290
rect 5347 3236 5353 3238
rect 5409 3236 5433 3238
rect 5489 3236 5513 3238
rect 5569 3236 5593 3238
rect 5649 3236 5655 3238
rect 5347 3227 5655 3236
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5736 2446 5764 4014
rect 5828 3194 5856 5510
rect 5920 5166 5948 6802
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 6842 6556 7150 6565
rect 6842 6554 6848 6556
rect 6904 6554 6928 6556
rect 6984 6554 7008 6556
rect 7064 6554 7088 6556
rect 7144 6554 7150 6556
rect 6904 6502 6906 6554
rect 7086 6502 7088 6554
rect 6842 6500 6848 6502
rect 6904 6500 6928 6502
rect 6984 6500 7008 6502
rect 7064 6500 7088 6502
rect 7144 6500 7150 6502
rect 6842 6491 7150 6500
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5920 2650 5948 5102
rect 6012 4826 6040 6190
rect 6182 6012 6490 6021
rect 6182 6010 6188 6012
rect 6244 6010 6268 6012
rect 6324 6010 6348 6012
rect 6404 6010 6428 6012
rect 6484 6010 6490 6012
rect 6244 5958 6246 6010
rect 6426 5958 6428 6010
rect 6182 5956 6188 5958
rect 6244 5956 6268 5958
rect 6324 5956 6348 5958
rect 6404 5956 6428 5958
rect 6484 5956 6490 5958
rect 6182 5947 6490 5956
rect 7300 5545 7328 6734
rect 7286 5536 7342 5545
rect 6842 5468 7150 5477
rect 7286 5471 7342 5480
rect 6842 5466 6848 5468
rect 6904 5466 6928 5468
rect 6984 5466 7008 5468
rect 7064 5466 7088 5468
rect 7144 5466 7150 5468
rect 6904 5414 6906 5466
rect 7086 5414 7088 5466
rect 6842 5412 6848 5414
rect 6904 5412 6928 5414
rect 6984 5412 7008 5414
rect 7064 5412 7088 5414
rect 7144 5412 7150 5414
rect 6842 5403 7150 5412
rect 6182 4924 6490 4933
rect 6182 4922 6188 4924
rect 6244 4922 6268 4924
rect 6324 4922 6348 4924
rect 6404 4922 6428 4924
rect 6484 4922 6490 4924
rect 6244 4870 6246 4922
rect 6426 4870 6428 4922
rect 6182 4868 6188 4870
rect 6244 4868 6268 4870
rect 6324 4868 6348 4870
rect 6404 4868 6428 4870
rect 6484 4868 6490 4870
rect 6182 4859 6490 4868
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6842 4380 7150 4389
rect 6842 4378 6848 4380
rect 6904 4378 6928 4380
rect 6984 4378 7008 4380
rect 7064 4378 7088 4380
rect 7144 4378 7150 4380
rect 6904 4326 6906 4378
rect 7086 4326 7088 4378
rect 6842 4324 6848 4326
rect 6904 4324 6928 4326
rect 6984 4324 7008 4326
rect 7064 4324 7088 4326
rect 7144 4324 7150 4326
rect 6842 4315 7150 4324
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6182 3836 6490 3845
rect 6182 3834 6188 3836
rect 6244 3834 6268 3836
rect 6324 3834 6348 3836
rect 6404 3834 6428 3836
rect 6484 3834 6490 3836
rect 6244 3782 6246 3834
rect 6426 3782 6428 3834
rect 6182 3780 6188 3782
rect 6244 3780 6268 3782
rect 6324 3780 6348 3782
rect 6404 3780 6428 3782
rect 6484 3780 6490 3782
rect 6182 3771 6490 3780
rect 6564 3738 6592 4014
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 3058 6040 3334
rect 6842 3292 7150 3301
rect 6842 3290 6848 3292
rect 6904 3290 6928 3292
rect 6984 3290 7008 3292
rect 7064 3290 7088 3292
rect 7144 3290 7150 3292
rect 6904 3238 6906 3290
rect 7086 3238 7088 3290
rect 6842 3236 6848 3238
rect 6904 3236 6928 3238
rect 6984 3236 7008 3238
rect 7064 3236 7088 3238
rect 7144 3236 7150 3238
rect 6842 3227 7150 3236
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6182 2748 6490 2757
rect 6182 2746 6188 2748
rect 6244 2746 6268 2748
rect 6324 2746 6348 2748
rect 6404 2746 6428 2748
rect 6484 2746 6490 2748
rect 6244 2694 6246 2746
rect 6426 2694 6428 2746
rect 6182 2692 6188 2694
rect 6244 2692 6268 2694
rect 6324 2692 6348 2694
rect 6404 2692 6428 2694
rect 6484 2692 6490 2694
rect 6182 2683 6490 2692
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 32 800 60 2246
rect 2357 2204 2665 2213
rect 2357 2202 2363 2204
rect 2419 2202 2443 2204
rect 2499 2202 2523 2204
rect 2579 2202 2603 2204
rect 2659 2202 2665 2204
rect 2419 2150 2421 2202
rect 2601 2150 2603 2202
rect 2357 2148 2363 2150
rect 2419 2148 2443 2150
rect 2499 2148 2523 2150
rect 2579 2148 2603 2150
rect 2659 2148 2665 2150
rect 2357 2139 2665 2148
rect 3252 800 3280 2246
rect 3852 2204 4160 2213
rect 3852 2202 3858 2204
rect 3914 2202 3938 2204
rect 3994 2202 4018 2204
rect 4074 2202 4098 2204
rect 4154 2202 4160 2204
rect 3914 2150 3916 2202
rect 4096 2150 4098 2202
rect 3852 2148 3858 2150
rect 3914 2148 3938 2150
rect 3994 2148 4018 2150
rect 4074 2148 4098 2150
rect 4154 2148 4160 2150
rect 3852 2139 4160 2148
rect 5347 2204 5655 2213
rect 5347 2202 5353 2204
rect 5409 2202 5433 2204
rect 5489 2202 5513 2204
rect 5569 2202 5593 2204
rect 5649 2202 5655 2204
rect 5409 2150 5411 2202
rect 5591 2150 5593 2202
rect 5347 2148 5353 2150
rect 5409 2148 5433 2150
rect 5489 2148 5513 2150
rect 5569 2148 5593 2150
rect 5649 2148 5655 2150
rect 5347 2139 5655 2148
rect 6472 800 6500 2246
rect 6842 2204 7150 2213
rect 6842 2202 6848 2204
rect 6904 2202 6928 2204
rect 6984 2202 7008 2204
rect 7064 2202 7088 2204
rect 7144 2202 7150 2204
rect 6904 2150 6906 2202
rect 7086 2150 7088 2202
rect 6842 2148 6848 2150
rect 6904 2148 6928 2150
rect 6984 2148 7008 2150
rect 7064 2148 7088 2150
rect 7144 2148 7150 2150
rect 6842 2139 7150 2148
rect 7300 1465 7328 2518
rect 7286 1456 7342 1465
rect 7286 1391 7342 1400
rect 18 0 74 800
rect 3238 0 3294 800
rect 6458 0 6514 800
<< via2 >>
rect 938 10240 994 10296
rect 1703 8186 1759 8188
rect 1783 8186 1839 8188
rect 1863 8186 1919 8188
rect 1943 8186 1999 8188
rect 1703 8134 1749 8186
rect 1749 8134 1759 8186
rect 1783 8134 1813 8186
rect 1813 8134 1825 8186
rect 1825 8134 1839 8186
rect 1863 8134 1877 8186
rect 1877 8134 1889 8186
rect 1889 8134 1919 8186
rect 1943 8134 1953 8186
rect 1953 8134 1999 8186
rect 1703 8132 1759 8134
rect 1783 8132 1839 8134
rect 1863 8132 1919 8134
rect 1943 8132 1999 8134
rect 3198 8186 3254 8188
rect 3278 8186 3334 8188
rect 3358 8186 3414 8188
rect 3438 8186 3494 8188
rect 3198 8134 3244 8186
rect 3244 8134 3254 8186
rect 3278 8134 3308 8186
rect 3308 8134 3320 8186
rect 3320 8134 3334 8186
rect 3358 8134 3372 8186
rect 3372 8134 3384 8186
rect 3384 8134 3414 8186
rect 3438 8134 3448 8186
rect 3448 8134 3494 8186
rect 3198 8132 3254 8134
rect 3278 8132 3334 8134
rect 3358 8132 3414 8134
rect 3438 8132 3494 8134
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4933 8186 4989 8188
rect 4693 8134 4739 8186
rect 4739 8134 4749 8186
rect 4773 8134 4803 8186
rect 4803 8134 4815 8186
rect 4815 8134 4829 8186
rect 4853 8134 4867 8186
rect 4867 8134 4879 8186
rect 4879 8134 4909 8186
rect 4933 8134 4943 8186
rect 4943 8134 4989 8186
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4933 8132 4989 8134
rect 7286 8880 7342 8936
rect 6188 8186 6244 8188
rect 6268 8186 6324 8188
rect 6348 8186 6404 8188
rect 6428 8186 6484 8188
rect 6188 8134 6234 8186
rect 6234 8134 6244 8186
rect 6268 8134 6298 8186
rect 6298 8134 6310 8186
rect 6310 8134 6324 8186
rect 6348 8134 6362 8186
rect 6362 8134 6374 8186
rect 6374 8134 6404 8186
rect 6428 8134 6438 8186
rect 6438 8134 6484 8186
rect 6188 8132 6244 8134
rect 6268 8132 6324 8134
rect 6348 8132 6404 8134
rect 6428 8132 6484 8134
rect 2363 7642 2419 7644
rect 2443 7642 2499 7644
rect 2523 7642 2579 7644
rect 2603 7642 2659 7644
rect 2363 7590 2409 7642
rect 2409 7590 2419 7642
rect 2443 7590 2473 7642
rect 2473 7590 2485 7642
rect 2485 7590 2499 7642
rect 2523 7590 2537 7642
rect 2537 7590 2549 7642
rect 2549 7590 2579 7642
rect 2603 7590 2613 7642
rect 2613 7590 2659 7642
rect 2363 7588 2419 7590
rect 2443 7588 2499 7590
rect 2523 7588 2579 7590
rect 2603 7588 2659 7590
rect 1703 7098 1759 7100
rect 1783 7098 1839 7100
rect 1863 7098 1919 7100
rect 1943 7098 1999 7100
rect 1703 7046 1749 7098
rect 1749 7046 1759 7098
rect 1783 7046 1813 7098
rect 1813 7046 1825 7098
rect 1825 7046 1839 7098
rect 1863 7046 1877 7098
rect 1877 7046 1889 7098
rect 1889 7046 1919 7098
rect 1943 7046 1953 7098
rect 1953 7046 1999 7098
rect 1703 7044 1759 7046
rect 1783 7044 1839 7046
rect 1863 7044 1919 7046
rect 1943 7044 1999 7046
rect 938 6840 994 6896
rect 3858 7642 3914 7644
rect 3938 7642 3994 7644
rect 4018 7642 4074 7644
rect 4098 7642 4154 7644
rect 3858 7590 3904 7642
rect 3904 7590 3914 7642
rect 3938 7590 3968 7642
rect 3968 7590 3980 7642
rect 3980 7590 3994 7642
rect 4018 7590 4032 7642
rect 4032 7590 4044 7642
rect 4044 7590 4074 7642
rect 4098 7590 4108 7642
rect 4108 7590 4154 7642
rect 3858 7588 3914 7590
rect 3938 7588 3994 7590
rect 4018 7588 4074 7590
rect 4098 7588 4154 7590
rect 1703 6010 1759 6012
rect 1783 6010 1839 6012
rect 1863 6010 1919 6012
rect 1943 6010 1999 6012
rect 1703 5958 1749 6010
rect 1749 5958 1759 6010
rect 1783 5958 1813 6010
rect 1813 5958 1825 6010
rect 1825 5958 1839 6010
rect 1863 5958 1877 6010
rect 1877 5958 1889 6010
rect 1889 5958 1919 6010
rect 1943 5958 1953 6010
rect 1953 5958 1999 6010
rect 1703 5956 1759 5958
rect 1783 5956 1839 5958
rect 1863 5956 1919 5958
rect 1943 5956 1999 5958
rect 1703 4922 1759 4924
rect 1783 4922 1839 4924
rect 1863 4922 1919 4924
rect 1943 4922 1999 4924
rect 1703 4870 1749 4922
rect 1749 4870 1759 4922
rect 1783 4870 1813 4922
rect 1813 4870 1825 4922
rect 1825 4870 1839 4922
rect 1863 4870 1877 4922
rect 1877 4870 1889 4922
rect 1889 4870 1919 4922
rect 1943 4870 1953 4922
rect 1953 4870 1999 4922
rect 1703 4868 1759 4870
rect 1783 4868 1839 4870
rect 1863 4868 1919 4870
rect 1943 4868 1999 4870
rect 1703 3834 1759 3836
rect 1783 3834 1839 3836
rect 1863 3834 1919 3836
rect 1943 3834 1999 3836
rect 1703 3782 1749 3834
rect 1749 3782 1759 3834
rect 1783 3782 1813 3834
rect 1813 3782 1825 3834
rect 1825 3782 1839 3834
rect 1863 3782 1877 3834
rect 1877 3782 1889 3834
rect 1889 3782 1919 3834
rect 1943 3782 1953 3834
rect 1953 3782 1999 3834
rect 1703 3780 1759 3782
rect 1783 3780 1839 3782
rect 1863 3780 1919 3782
rect 1943 3780 1999 3782
rect 938 3440 994 3496
rect 2363 6554 2419 6556
rect 2443 6554 2499 6556
rect 2523 6554 2579 6556
rect 2603 6554 2659 6556
rect 2363 6502 2409 6554
rect 2409 6502 2419 6554
rect 2443 6502 2473 6554
rect 2473 6502 2485 6554
rect 2485 6502 2499 6554
rect 2523 6502 2537 6554
rect 2537 6502 2549 6554
rect 2549 6502 2579 6554
rect 2603 6502 2613 6554
rect 2613 6502 2659 6554
rect 2363 6500 2419 6502
rect 2443 6500 2499 6502
rect 2523 6500 2579 6502
rect 2603 6500 2659 6502
rect 2363 5466 2419 5468
rect 2443 5466 2499 5468
rect 2523 5466 2579 5468
rect 2603 5466 2659 5468
rect 2363 5414 2409 5466
rect 2409 5414 2419 5466
rect 2443 5414 2473 5466
rect 2473 5414 2485 5466
rect 2485 5414 2499 5466
rect 2523 5414 2537 5466
rect 2537 5414 2549 5466
rect 2549 5414 2579 5466
rect 2603 5414 2613 5466
rect 2613 5414 2659 5466
rect 2363 5412 2419 5414
rect 2443 5412 2499 5414
rect 2523 5412 2579 5414
rect 2603 5412 2659 5414
rect 2363 4378 2419 4380
rect 2443 4378 2499 4380
rect 2523 4378 2579 4380
rect 2603 4378 2659 4380
rect 2363 4326 2409 4378
rect 2409 4326 2419 4378
rect 2443 4326 2473 4378
rect 2473 4326 2485 4378
rect 2485 4326 2499 4378
rect 2523 4326 2537 4378
rect 2537 4326 2549 4378
rect 2549 4326 2579 4378
rect 2603 4326 2613 4378
rect 2613 4326 2659 4378
rect 2363 4324 2419 4326
rect 2443 4324 2499 4326
rect 2523 4324 2579 4326
rect 2603 4324 2659 4326
rect 2363 3290 2419 3292
rect 2443 3290 2499 3292
rect 2523 3290 2579 3292
rect 2603 3290 2659 3292
rect 2363 3238 2409 3290
rect 2409 3238 2419 3290
rect 2443 3238 2473 3290
rect 2473 3238 2485 3290
rect 2485 3238 2499 3290
rect 2523 3238 2537 3290
rect 2537 3238 2549 3290
rect 2549 3238 2579 3290
rect 2603 3238 2613 3290
rect 2613 3238 2659 3290
rect 2363 3236 2419 3238
rect 2443 3236 2499 3238
rect 2523 3236 2579 3238
rect 2603 3236 2659 3238
rect 1703 2746 1759 2748
rect 1783 2746 1839 2748
rect 1863 2746 1919 2748
rect 1943 2746 1999 2748
rect 1703 2694 1749 2746
rect 1749 2694 1759 2746
rect 1783 2694 1813 2746
rect 1813 2694 1825 2746
rect 1825 2694 1839 2746
rect 1863 2694 1877 2746
rect 1877 2694 1889 2746
rect 1889 2694 1919 2746
rect 1943 2694 1953 2746
rect 1953 2694 1999 2746
rect 1703 2692 1759 2694
rect 1783 2692 1839 2694
rect 1863 2692 1919 2694
rect 1943 2692 1999 2694
rect 3198 7098 3254 7100
rect 3278 7098 3334 7100
rect 3358 7098 3414 7100
rect 3438 7098 3494 7100
rect 3198 7046 3244 7098
rect 3244 7046 3254 7098
rect 3278 7046 3308 7098
rect 3308 7046 3320 7098
rect 3320 7046 3334 7098
rect 3358 7046 3372 7098
rect 3372 7046 3384 7098
rect 3384 7046 3414 7098
rect 3438 7046 3448 7098
rect 3448 7046 3494 7098
rect 3198 7044 3254 7046
rect 3278 7044 3334 7046
rect 3358 7044 3414 7046
rect 3438 7044 3494 7046
rect 3858 6554 3914 6556
rect 3938 6554 3994 6556
rect 4018 6554 4074 6556
rect 4098 6554 4154 6556
rect 3858 6502 3904 6554
rect 3904 6502 3914 6554
rect 3938 6502 3968 6554
rect 3968 6502 3980 6554
rect 3980 6502 3994 6554
rect 4018 6502 4032 6554
rect 4032 6502 4044 6554
rect 4044 6502 4074 6554
rect 4098 6502 4108 6554
rect 4108 6502 4154 6554
rect 3858 6500 3914 6502
rect 3938 6500 3994 6502
rect 4018 6500 4074 6502
rect 4098 6500 4154 6502
rect 3198 6010 3254 6012
rect 3278 6010 3334 6012
rect 3358 6010 3414 6012
rect 3438 6010 3494 6012
rect 3198 5958 3244 6010
rect 3244 5958 3254 6010
rect 3278 5958 3308 6010
rect 3308 5958 3320 6010
rect 3320 5958 3334 6010
rect 3358 5958 3372 6010
rect 3372 5958 3384 6010
rect 3384 5958 3414 6010
rect 3438 5958 3448 6010
rect 3448 5958 3494 6010
rect 3198 5956 3254 5958
rect 3278 5956 3334 5958
rect 3358 5956 3414 5958
rect 3438 5956 3494 5958
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4933 7098 4989 7100
rect 4693 7046 4739 7098
rect 4739 7046 4749 7098
rect 4773 7046 4803 7098
rect 4803 7046 4815 7098
rect 4815 7046 4829 7098
rect 4853 7046 4867 7098
rect 4867 7046 4879 7098
rect 4879 7046 4909 7098
rect 4933 7046 4943 7098
rect 4943 7046 4989 7098
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4933 7044 4989 7046
rect 3858 5466 3914 5468
rect 3938 5466 3994 5468
rect 4018 5466 4074 5468
rect 4098 5466 4154 5468
rect 3858 5414 3904 5466
rect 3904 5414 3914 5466
rect 3938 5414 3968 5466
rect 3968 5414 3980 5466
rect 3980 5414 3994 5466
rect 4018 5414 4032 5466
rect 4032 5414 4044 5466
rect 4044 5414 4074 5466
rect 4098 5414 4108 5466
rect 4108 5414 4154 5466
rect 3858 5412 3914 5414
rect 3938 5412 3994 5414
rect 4018 5412 4074 5414
rect 4098 5412 4154 5414
rect 3198 4922 3254 4924
rect 3278 4922 3334 4924
rect 3358 4922 3414 4924
rect 3438 4922 3494 4924
rect 3198 4870 3244 4922
rect 3244 4870 3254 4922
rect 3278 4870 3308 4922
rect 3308 4870 3320 4922
rect 3320 4870 3334 4922
rect 3358 4870 3372 4922
rect 3372 4870 3384 4922
rect 3384 4870 3414 4922
rect 3438 4870 3448 4922
rect 3448 4870 3494 4922
rect 3198 4868 3254 4870
rect 3278 4868 3334 4870
rect 3358 4868 3414 4870
rect 3438 4868 3494 4870
rect 3198 3834 3254 3836
rect 3278 3834 3334 3836
rect 3358 3834 3414 3836
rect 3438 3834 3494 3836
rect 3198 3782 3244 3834
rect 3244 3782 3254 3834
rect 3278 3782 3308 3834
rect 3308 3782 3320 3834
rect 3320 3782 3334 3834
rect 3358 3782 3372 3834
rect 3372 3782 3384 3834
rect 3384 3782 3414 3834
rect 3438 3782 3448 3834
rect 3448 3782 3494 3834
rect 3198 3780 3254 3782
rect 3278 3780 3334 3782
rect 3358 3780 3414 3782
rect 3438 3780 3494 3782
rect 3198 2746 3254 2748
rect 3278 2746 3334 2748
rect 3358 2746 3414 2748
rect 3438 2746 3494 2748
rect 3198 2694 3244 2746
rect 3244 2694 3254 2746
rect 3278 2694 3308 2746
rect 3308 2694 3320 2746
rect 3320 2694 3334 2746
rect 3358 2694 3372 2746
rect 3372 2694 3384 2746
rect 3384 2694 3414 2746
rect 3438 2694 3448 2746
rect 3448 2694 3494 2746
rect 3198 2692 3254 2694
rect 3278 2692 3334 2694
rect 3358 2692 3414 2694
rect 3438 2692 3494 2694
rect 3858 4378 3914 4380
rect 3938 4378 3994 4380
rect 4018 4378 4074 4380
rect 4098 4378 4154 4380
rect 3858 4326 3904 4378
rect 3904 4326 3914 4378
rect 3938 4326 3968 4378
rect 3968 4326 3980 4378
rect 3980 4326 3994 4378
rect 4018 4326 4032 4378
rect 4032 4326 4044 4378
rect 4044 4326 4074 4378
rect 4098 4326 4108 4378
rect 4108 4326 4154 4378
rect 3858 4324 3914 4326
rect 3938 4324 3994 4326
rect 4018 4324 4074 4326
rect 4098 4324 4154 4326
rect 3858 3290 3914 3292
rect 3938 3290 3994 3292
rect 4018 3290 4074 3292
rect 4098 3290 4154 3292
rect 3858 3238 3904 3290
rect 3904 3238 3914 3290
rect 3938 3238 3968 3290
rect 3968 3238 3980 3290
rect 3980 3238 3994 3290
rect 4018 3238 4032 3290
rect 4032 3238 4044 3290
rect 4044 3238 4074 3290
rect 4098 3238 4108 3290
rect 4108 3238 4154 3290
rect 3858 3236 3914 3238
rect 3938 3236 3994 3238
rect 4018 3236 4074 3238
rect 4098 3236 4154 3238
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4933 6010 4989 6012
rect 4693 5958 4739 6010
rect 4739 5958 4749 6010
rect 4773 5958 4803 6010
rect 4803 5958 4815 6010
rect 4815 5958 4829 6010
rect 4853 5958 4867 6010
rect 4867 5958 4879 6010
rect 4879 5958 4909 6010
rect 4933 5958 4943 6010
rect 4943 5958 4989 6010
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4933 5956 4989 5958
rect 5353 7642 5409 7644
rect 5433 7642 5489 7644
rect 5513 7642 5569 7644
rect 5593 7642 5649 7644
rect 5353 7590 5399 7642
rect 5399 7590 5409 7642
rect 5433 7590 5463 7642
rect 5463 7590 5475 7642
rect 5475 7590 5489 7642
rect 5513 7590 5527 7642
rect 5527 7590 5539 7642
rect 5539 7590 5569 7642
rect 5593 7590 5603 7642
rect 5603 7590 5649 7642
rect 5353 7588 5409 7590
rect 5433 7588 5489 7590
rect 5513 7588 5569 7590
rect 5593 7588 5649 7590
rect 6848 7642 6904 7644
rect 6928 7642 6984 7644
rect 7008 7642 7064 7644
rect 7088 7642 7144 7644
rect 6848 7590 6894 7642
rect 6894 7590 6904 7642
rect 6928 7590 6958 7642
rect 6958 7590 6970 7642
rect 6970 7590 6984 7642
rect 7008 7590 7022 7642
rect 7022 7590 7034 7642
rect 7034 7590 7064 7642
rect 7088 7590 7098 7642
rect 7098 7590 7144 7642
rect 6848 7588 6904 7590
rect 6928 7588 6984 7590
rect 7008 7588 7064 7590
rect 7088 7588 7144 7590
rect 6188 7098 6244 7100
rect 6268 7098 6324 7100
rect 6348 7098 6404 7100
rect 6428 7098 6484 7100
rect 6188 7046 6234 7098
rect 6234 7046 6244 7098
rect 6268 7046 6298 7098
rect 6298 7046 6310 7098
rect 6310 7046 6324 7098
rect 6348 7046 6362 7098
rect 6362 7046 6374 7098
rect 6374 7046 6404 7098
rect 6428 7046 6438 7098
rect 6438 7046 6484 7098
rect 6188 7044 6244 7046
rect 6268 7044 6324 7046
rect 6348 7044 6404 7046
rect 6428 7044 6484 7046
rect 5353 6554 5409 6556
rect 5433 6554 5489 6556
rect 5513 6554 5569 6556
rect 5593 6554 5649 6556
rect 5353 6502 5399 6554
rect 5399 6502 5409 6554
rect 5433 6502 5463 6554
rect 5463 6502 5475 6554
rect 5475 6502 5489 6554
rect 5513 6502 5527 6554
rect 5527 6502 5539 6554
rect 5539 6502 5569 6554
rect 5593 6502 5603 6554
rect 5603 6502 5649 6554
rect 5353 6500 5409 6502
rect 5433 6500 5489 6502
rect 5513 6500 5569 6502
rect 5593 6500 5649 6502
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4933 4922 4989 4924
rect 4693 4870 4739 4922
rect 4739 4870 4749 4922
rect 4773 4870 4803 4922
rect 4803 4870 4815 4922
rect 4815 4870 4829 4922
rect 4853 4870 4867 4922
rect 4867 4870 4879 4922
rect 4879 4870 4909 4922
rect 4933 4870 4943 4922
rect 4943 4870 4989 4922
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4933 4868 4989 4870
rect 5353 5466 5409 5468
rect 5433 5466 5489 5468
rect 5513 5466 5569 5468
rect 5593 5466 5649 5468
rect 5353 5414 5399 5466
rect 5399 5414 5409 5466
rect 5433 5414 5463 5466
rect 5463 5414 5475 5466
rect 5475 5414 5489 5466
rect 5513 5414 5527 5466
rect 5527 5414 5539 5466
rect 5539 5414 5569 5466
rect 5593 5414 5603 5466
rect 5603 5414 5649 5466
rect 5353 5412 5409 5414
rect 5433 5412 5489 5414
rect 5513 5412 5569 5414
rect 5593 5412 5649 5414
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4933 3834 4989 3836
rect 4693 3782 4739 3834
rect 4739 3782 4749 3834
rect 4773 3782 4803 3834
rect 4803 3782 4815 3834
rect 4815 3782 4829 3834
rect 4853 3782 4867 3834
rect 4867 3782 4879 3834
rect 4879 3782 4909 3834
rect 4933 3782 4943 3834
rect 4943 3782 4989 3834
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4933 3780 4989 3782
rect 5353 4378 5409 4380
rect 5433 4378 5489 4380
rect 5513 4378 5569 4380
rect 5593 4378 5649 4380
rect 5353 4326 5399 4378
rect 5399 4326 5409 4378
rect 5433 4326 5463 4378
rect 5463 4326 5475 4378
rect 5475 4326 5489 4378
rect 5513 4326 5527 4378
rect 5527 4326 5539 4378
rect 5539 4326 5569 4378
rect 5593 4326 5603 4378
rect 5603 4326 5649 4378
rect 5353 4324 5409 4326
rect 5433 4324 5489 4326
rect 5513 4324 5569 4326
rect 5593 4324 5649 4326
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4933 2746 4989 2748
rect 4693 2694 4739 2746
rect 4739 2694 4749 2746
rect 4773 2694 4803 2746
rect 4803 2694 4815 2746
rect 4815 2694 4829 2746
rect 4853 2694 4867 2746
rect 4867 2694 4879 2746
rect 4879 2694 4909 2746
rect 4933 2694 4943 2746
rect 4943 2694 4989 2746
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 4933 2692 4989 2694
rect 5353 3290 5409 3292
rect 5433 3290 5489 3292
rect 5513 3290 5569 3292
rect 5593 3290 5649 3292
rect 5353 3238 5399 3290
rect 5399 3238 5409 3290
rect 5433 3238 5463 3290
rect 5463 3238 5475 3290
rect 5475 3238 5489 3290
rect 5513 3238 5527 3290
rect 5527 3238 5539 3290
rect 5539 3238 5569 3290
rect 5593 3238 5603 3290
rect 5603 3238 5649 3290
rect 5353 3236 5409 3238
rect 5433 3236 5489 3238
rect 5513 3236 5569 3238
rect 5593 3236 5649 3238
rect 6848 6554 6904 6556
rect 6928 6554 6984 6556
rect 7008 6554 7064 6556
rect 7088 6554 7144 6556
rect 6848 6502 6894 6554
rect 6894 6502 6904 6554
rect 6928 6502 6958 6554
rect 6958 6502 6970 6554
rect 6970 6502 6984 6554
rect 7008 6502 7022 6554
rect 7022 6502 7034 6554
rect 7034 6502 7064 6554
rect 7088 6502 7098 6554
rect 7098 6502 7144 6554
rect 6848 6500 6904 6502
rect 6928 6500 6984 6502
rect 7008 6500 7064 6502
rect 7088 6500 7144 6502
rect 6188 6010 6244 6012
rect 6268 6010 6324 6012
rect 6348 6010 6404 6012
rect 6428 6010 6484 6012
rect 6188 5958 6234 6010
rect 6234 5958 6244 6010
rect 6268 5958 6298 6010
rect 6298 5958 6310 6010
rect 6310 5958 6324 6010
rect 6348 5958 6362 6010
rect 6362 5958 6374 6010
rect 6374 5958 6404 6010
rect 6428 5958 6438 6010
rect 6438 5958 6484 6010
rect 6188 5956 6244 5958
rect 6268 5956 6324 5958
rect 6348 5956 6404 5958
rect 6428 5956 6484 5958
rect 7286 5480 7342 5536
rect 6848 5466 6904 5468
rect 6928 5466 6984 5468
rect 7008 5466 7064 5468
rect 7088 5466 7144 5468
rect 6848 5414 6894 5466
rect 6894 5414 6904 5466
rect 6928 5414 6958 5466
rect 6958 5414 6970 5466
rect 6970 5414 6984 5466
rect 7008 5414 7022 5466
rect 7022 5414 7034 5466
rect 7034 5414 7064 5466
rect 7088 5414 7098 5466
rect 7098 5414 7144 5466
rect 6848 5412 6904 5414
rect 6928 5412 6984 5414
rect 7008 5412 7064 5414
rect 7088 5412 7144 5414
rect 6188 4922 6244 4924
rect 6268 4922 6324 4924
rect 6348 4922 6404 4924
rect 6428 4922 6484 4924
rect 6188 4870 6234 4922
rect 6234 4870 6244 4922
rect 6268 4870 6298 4922
rect 6298 4870 6310 4922
rect 6310 4870 6324 4922
rect 6348 4870 6362 4922
rect 6362 4870 6374 4922
rect 6374 4870 6404 4922
rect 6428 4870 6438 4922
rect 6438 4870 6484 4922
rect 6188 4868 6244 4870
rect 6268 4868 6324 4870
rect 6348 4868 6404 4870
rect 6428 4868 6484 4870
rect 6848 4378 6904 4380
rect 6928 4378 6984 4380
rect 7008 4378 7064 4380
rect 7088 4378 7144 4380
rect 6848 4326 6894 4378
rect 6894 4326 6904 4378
rect 6928 4326 6958 4378
rect 6958 4326 6970 4378
rect 6970 4326 6984 4378
rect 7008 4326 7022 4378
rect 7022 4326 7034 4378
rect 7034 4326 7064 4378
rect 7088 4326 7098 4378
rect 7098 4326 7144 4378
rect 6848 4324 6904 4326
rect 6928 4324 6984 4326
rect 7008 4324 7064 4326
rect 7088 4324 7144 4326
rect 6188 3834 6244 3836
rect 6268 3834 6324 3836
rect 6348 3834 6404 3836
rect 6428 3834 6484 3836
rect 6188 3782 6234 3834
rect 6234 3782 6244 3834
rect 6268 3782 6298 3834
rect 6298 3782 6310 3834
rect 6310 3782 6324 3834
rect 6348 3782 6362 3834
rect 6362 3782 6374 3834
rect 6374 3782 6404 3834
rect 6428 3782 6438 3834
rect 6438 3782 6484 3834
rect 6188 3780 6244 3782
rect 6268 3780 6324 3782
rect 6348 3780 6404 3782
rect 6428 3780 6484 3782
rect 6848 3290 6904 3292
rect 6928 3290 6984 3292
rect 7008 3290 7064 3292
rect 7088 3290 7144 3292
rect 6848 3238 6894 3290
rect 6894 3238 6904 3290
rect 6928 3238 6958 3290
rect 6958 3238 6970 3290
rect 6970 3238 6984 3290
rect 7008 3238 7022 3290
rect 7022 3238 7034 3290
rect 7034 3238 7064 3290
rect 7088 3238 7098 3290
rect 7098 3238 7144 3290
rect 6848 3236 6904 3238
rect 6928 3236 6984 3238
rect 7008 3236 7064 3238
rect 7088 3236 7144 3238
rect 6188 2746 6244 2748
rect 6268 2746 6324 2748
rect 6348 2746 6404 2748
rect 6428 2746 6484 2748
rect 6188 2694 6234 2746
rect 6234 2694 6244 2746
rect 6268 2694 6298 2746
rect 6298 2694 6310 2746
rect 6310 2694 6324 2746
rect 6348 2694 6362 2746
rect 6362 2694 6374 2746
rect 6374 2694 6404 2746
rect 6428 2694 6438 2746
rect 6438 2694 6484 2746
rect 6188 2692 6244 2694
rect 6268 2692 6324 2694
rect 6348 2692 6404 2694
rect 6428 2692 6484 2694
rect 2363 2202 2419 2204
rect 2443 2202 2499 2204
rect 2523 2202 2579 2204
rect 2603 2202 2659 2204
rect 2363 2150 2409 2202
rect 2409 2150 2419 2202
rect 2443 2150 2473 2202
rect 2473 2150 2485 2202
rect 2485 2150 2499 2202
rect 2523 2150 2537 2202
rect 2537 2150 2549 2202
rect 2549 2150 2579 2202
rect 2603 2150 2613 2202
rect 2613 2150 2659 2202
rect 2363 2148 2419 2150
rect 2443 2148 2499 2150
rect 2523 2148 2579 2150
rect 2603 2148 2659 2150
rect 3858 2202 3914 2204
rect 3938 2202 3994 2204
rect 4018 2202 4074 2204
rect 4098 2202 4154 2204
rect 3858 2150 3904 2202
rect 3904 2150 3914 2202
rect 3938 2150 3968 2202
rect 3968 2150 3980 2202
rect 3980 2150 3994 2202
rect 4018 2150 4032 2202
rect 4032 2150 4044 2202
rect 4044 2150 4074 2202
rect 4098 2150 4108 2202
rect 4108 2150 4154 2202
rect 3858 2148 3914 2150
rect 3938 2148 3994 2150
rect 4018 2148 4074 2150
rect 4098 2148 4154 2150
rect 5353 2202 5409 2204
rect 5433 2202 5489 2204
rect 5513 2202 5569 2204
rect 5593 2202 5649 2204
rect 5353 2150 5399 2202
rect 5399 2150 5409 2202
rect 5433 2150 5463 2202
rect 5463 2150 5475 2202
rect 5475 2150 5489 2202
rect 5513 2150 5527 2202
rect 5527 2150 5539 2202
rect 5539 2150 5569 2202
rect 5593 2150 5603 2202
rect 5603 2150 5649 2202
rect 5353 2148 5409 2150
rect 5433 2148 5489 2150
rect 5513 2148 5569 2150
rect 5593 2148 5649 2150
rect 6848 2202 6904 2204
rect 6928 2202 6984 2204
rect 7008 2202 7064 2204
rect 7088 2202 7144 2204
rect 6848 2150 6894 2202
rect 6894 2150 6904 2202
rect 6928 2150 6958 2202
rect 6958 2150 6970 2202
rect 6970 2150 6984 2202
rect 7008 2150 7022 2202
rect 7022 2150 7034 2202
rect 7034 2150 7064 2202
rect 7088 2150 7098 2202
rect 7098 2150 7144 2202
rect 6848 2148 6904 2150
rect 6928 2148 6984 2150
rect 7008 2148 7064 2150
rect 7088 2148 7144 2150
rect 7286 1400 7342 1456
<< metal3 >>
rect 0 10298 800 10328
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 7281 8938 7347 8941
rect 7458 8938 8258 8968
rect 7281 8936 8258 8938
rect 7281 8880 7286 8936
rect 7342 8880 8258 8936
rect 7281 8878 8258 8880
rect 7281 8875 7347 8878
rect 7458 8848 8258 8878
rect 1693 8192 2009 8193
rect 1693 8128 1699 8192
rect 1763 8128 1779 8192
rect 1843 8128 1859 8192
rect 1923 8128 1939 8192
rect 2003 8128 2009 8192
rect 1693 8127 2009 8128
rect 3188 8192 3504 8193
rect 3188 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3434 8192
rect 3498 8128 3504 8192
rect 3188 8127 3504 8128
rect 4683 8192 4999 8193
rect 4683 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4929 8192
rect 4993 8128 4999 8192
rect 4683 8127 4999 8128
rect 6178 8192 6494 8193
rect 6178 8128 6184 8192
rect 6248 8128 6264 8192
rect 6328 8128 6344 8192
rect 6408 8128 6424 8192
rect 6488 8128 6494 8192
rect 6178 8127 6494 8128
rect 2353 7648 2669 7649
rect 2353 7584 2359 7648
rect 2423 7584 2439 7648
rect 2503 7584 2519 7648
rect 2583 7584 2599 7648
rect 2663 7584 2669 7648
rect 2353 7583 2669 7584
rect 3848 7648 4164 7649
rect 3848 7584 3854 7648
rect 3918 7584 3934 7648
rect 3998 7584 4014 7648
rect 4078 7584 4094 7648
rect 4158 7584 4164 7648
rect 3848 7583 4164 7584
rect 5343 7648 5659 7649
rect 5343 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5589 7648
rect 5653 7584 5659 7648
rect 5343 7583 5659 7584
rect 6838 7648 7154 7649
rect 6838 7584 6844 7648
rect 6908 7584 6924 7648
rect 6988 7584 7004 7648
rect 7068 7584 7084 7648
rect 7148 7584 7154 7648
rect 6838 7583 7154 7584
rect 1693 7104 2009 7105
rect 1693 7040 1699 7104
rect 1763 7040 1779 7104
rect 1843 7040 1859 7104
rect 1923 7040 1939 7104
rect 2003 7040 2009 7104
rect 1693 7039 2009 7040
rect 3188 7104 3504 7105
rect 3188 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3434 7104
rect 3498 7040 3504 7104
rect 3188 7039 3504 7040
rect 4683 7104 4999 7105
rect 4683 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4929 7104
rect 4993 7040 4999 7104
rect 4683 7039 4999 7040
rect 6178 7104 6494 7105
rect 6178 7040 6184 7104
rect 6248 7040 6264 7104
rect 6328 7040 6344 7104
rect 6408 7040 6424 7104
rect 6488 7040 6494 7104
rect 6178 7039 6494 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 2353 6560 2669 6561
rect 2353 6496 2359 6560
rect 2423 6496 2439 6560
rect 2503 6496 2519 6560
rect 2583 6496 2599 6560
rect 2663 6496 2669 6560
rect 2353 6495 2669 6496
rect 3848 6560 4164 6561
rect 3848 6496 3854 6560
rect 3918 6496 3934 6560
rect 3998 6496 4014 6560
rect 4078 6496 4094 6560
rect 4158 6496 4164 6560
rect 3848 6495 4164 6496
rect 5343 6560 5659 6561
rect 5343 6496 5349 6560
rect 5413 6496 5429 6560
rect 5493 6496 5509 6560
rect 5573 6496 5589 6560
rect 5653 6496 5659 6560
rect 5343 6495 5659 6496
rect 6838 6560 7154 6561
rect 6838 6496 6844 6560
rect 6908 6496 6924 6560
rect 6988 6496 7004 6560
rect 7068 6496 7084 6560
rect 7148 6496 7154 6560
rect 6838 6495 7154 6496
rect 1693 6016 2009 6017
rect 1693 5952 1699 6016
rect 1763 5952 1779 6016
rect 1843 5952 1859 6016
rect 1923 5952 1939 6016
rect 2003 5952 2009 6016
rect 1693 5951 2009 5952
rect 3188 6016 3504 6017
rect 3188 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3434 6016
rect 3498 5952 3504 6016
rect 3188 5951 3504 5952
rect 4683 6016 4999 6017
rect 4683 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4929 6016
rect 4993 5952 4999 6016
rect 4683 5951 4999 5952
rect 6178 6016 6494 6017
rect 6178 5952 6184 6016
rect 6248 5952 6264 6016
rect 6328 5952 6344 6016
rect 6408 5952 6424 6016
rect 6488 5952 6494 6016
rect 6178 5951 6494 5952
rect 7281 5538 7347 5541
rect 7458 5538 8258 5568
rect 7281 5536 8258 5538
rect 7281 5480 7286 5536
rect 7342 5480 8258 5536
rect 7281 5478 8258 5480
rect 7281 5475 7347 5478
rect 2353 5472 2669 5473
rect 2353 5408 2359 5472
rect 2423 5408 2439 5472
rect 2503 5408 2519 5472
rect 2583 5408 2599 5472
rect 2663 5408 2669 5472
rect 2353 5407 2669 5408
rect 3848 5472 4164 5473
rect 3848 5408 3854 5472
rect 3918 5408 3934 5472
rect 3998 5408 4014 5472
rect 4078 5408 4094 5472
rect 4158 5408 4164 5472
rect 3848 5407 4164 5408
rect 5343 5472 5659 5473
rect 5343 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5589 5472
rect 5653 5408 5659 5472
rect 5343 5407 5659 5408
rect 6838 5472 7154 5473
rect 6838 5408 6844 5472
rect 6908 5408 6924 5472
rect 6988 5408 7004 5472
rect 7068 5408 7084 5472
rect 7148 5408 7154 5472
rect 7458 5448 8258 5478
rect 6838 5407 7154 5408
rect 1693 4928 2009 4929
rect 1693 4864 1699 4928
rect 1763 4864 1779 4928
rect 1843 4864 1859 4928
rect 1923 4864 1939 4928
rect 2003 4864 2009 4928
rect 1693 4863 2009 4864
rect 3188 4928 3504 4929
rect 3188 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3434 4928
rect 3498 4864 3504 4928
rect 3188 4863 3504 4864
rect 4683 4928 4999 4929
rect 4683 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4929 4928
rect 4993 4864 4999 4928
rect 4683 4863 4999 4864
rect 6178 4928 6494 4929
rect 6178 4864 6184 4928
rect 6248 4864 6264 4928
rect 6328 4864 6344 4928
rect 6408 4864 6424 4928
rect 6488 4864 6494 4928
rect 6178 4863 6494 4864
rect 2353 4384 2669 4385
rect 2353 4320 2359 4384
rect 2423 4320 2439 4384
rect 2503 4320 2519 4384
rect 2583 4320 2599 4384
rect 2663 4320 2669 4384
rect 2353 4319 2669 4320
rect 3848 4384 4164 4385
rect 3848 4320 3854 4384
rect 3918 4320 3934 4384
rect 3998 4320 4014 4384
rect 4078 4320 4094 4384
rect 4158 4320 4164 4384
rect 3848 4319 4164 4320
rect 5343 4384 5659 4385
rect 5343 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5589 4384
rect 5653 4320 5659 4384
rect 5343 4319 5659 4320
rect 6838 4384 7154 4385
rect 6838 4320 6844 4384
rect 6908 4320 6924 4384
rect 6988 4320 7004 4384
rect 7068 4320 7084 4384
rect 7148 4320 7154 4384
rect 6838 4319 7154 4320
rect 1693 3840 2009 3841
rect 1693 3776 1699 3840
rect 1763 3776 1779 3840
rect 1843 3776 1859 3840
rect 1923 3776 1939 3840
rect 2003 3776 2009 3840
rect 1693 3775 2009 3776
rect 3188 3840 3504 3841
rect 3188 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3434 3840
rect 3498 3776 3504 3840
rect 3188 3775 3504 3776
rect 4683 3840 4999 3841
rect 4683 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4929 3840
rect 4993 3776 4999 3840
rect 4683 3775 4999 3776
rect 6178 3840 6494 3841
rect 6178 3776 6184 3840
rect 6248 3776 6264 3840
rect 6328 3776 6344 3840
rect 6408 3776 6424 3840
rect 6488 3776 6494 3840
rect 6178 3775 6494 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 2353 3296 2669 3297
rect 2353 3232 2359 3296
rect 2423 3232 2439 3296
rect 2503 3232 2519 3296
rect 2583 3232 2599 3296
rect 2663 3232 2669 3296
rect 2353 3231 2669 3232
rect 3848 3296 4164 3297
rect 3848 3232 3854 3296
rect 3918 3232 3934 3296
rect 3998 3232 4014 3296
rect 4078 3232 4094 3296
rect 4158 3232 4164 3296
rect 3848 3231 4164 3232
rect 5343 3296 5659 3297
rect 5343 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5589 3296
rect 5653 3232 5659 3296
rect 5343 3231 5659 3232
rect 6838 3296 7154 3297
rect 6838 3232 6844 3296
rect 6908 3232 6924 3296
rect 6988 3232 7004 3296
rect 7068 3232 7084 3296
rect 7148 3232 7154 3296
rect 6838 3231 7154 3232
rect 1693 2752 2009 2753
rect 1693 2688 1699 2752
rect 1763 2688 1779 2752
rect 1843 2688 1859 2752
rect 1923 2688 1939 2752
rect 2003 2688 2009 2752
rect 1693 2687 2009 2688
rect 3188 2752 3504 2753
rect 3188 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3434 2752
rect 3498 2688 3504 2752
rect 3188 2687 3504 2688
rect 4683 2752 4999 2753
rect 4683 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4929 2752
rect 4993 2688 4999 2752
rect 4683 2687 4999 2688
rect 6178 2752 6494 2753
rect 6178 2688 6184 2752
rect 6248 2688 6264 2752
rect 6328 2688 6344 2752
rect 6408 2688 6424 2752
rect 6488 2688 6494 2752
rect 6178 2687 6494 2688
rect 2353 2208 2669 2209
rect 2353 2144 2359 2208
rect 2423 2144 2439 2208
rect 2503 2144 2519 2208
rect 2583 2144 2599 2208
rect 2663 2144 2669 2208
rect 2353 2143 2669 2144
rect 3848 2208 4164 2209
rect 3848 2144 3854 2208
rect 3918 2144 3934 2208
rect 3998 2144 4014 2208
rect 4078 2144 4094 2208
rect 4158 2144 4164 2208
rect 3848 2143 4164 2144
rect 5343 2208 5659 2209
rect 5343 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5589 2208
rect 5653 2144 5659 2208
rect 5343 2143 5659 2144
rect 6838 2208 7154 2209
rect 6838 2144 6844 2208
rect 6908 2144 6924 2208
rect 6988 2144 7004 2208
rect 7068 2144 7084 2208
rect 7148 2144 7154 2208
rect 6838 2143 7154 2144
rect 7281 1458 7347 1461
rect 7458 1458 8258 1488
rect 7281 1456 8258 1458
rect 7281 1400 7286 1456
rect 7342 1400 8258 1456
rect 7281 1398 8258 1400
rect 7281 1395 7347 1398
rect 7458 1368 8258 1398
<< via3 >>
rect 1699 8188 1763 8192
rect 1699 8132 1703 8188
rect 1703 8132 1759 8188
rect 1759 8132 1763 8188
rect 1699 8128 1763 8132
rect 1779 8188 1843 8192
rect 1779 8132 1783 8188
rect 1783 8132 1839 8188
rect 1839 8132 1843 8188
rect 1779 8128 1843 8132
rect 1859 8188 1923 8192
rect 1859 8132 1863 8188
rect 1863 8132 1919 8188
rect 1919 8132 1923 8188
rect 1859 8128 1923 8132
rect 1939 8188 2003 8192
rect 1939 8132 1943 8188
rect 1943 8132 1999 8188
rect 1999 8132 2003 8188
rect 1939 8128 2003 8132
rect 3194 8188 3258 8192
rect 3194 8132 3198 8188
rect 3198 8132 3254 8188
rect 3254 8132 3258 8188
rect 3194 8128 3258 8132
rect 3274 8188 3338 8192
rect 3274 8132 3278 8188
rect 3278 8132 3334 8188
rect 3334 8132 3338 8188
rect 3274 8128 3338 8132
rect 3354 8188 3418 8192
rect 3354 8132 3358 8188
rect 3358 8132 3414 8188
rect 3414 8132 3418 8188
rect 3354 8128 3418 8132
rect 3434 8188 3498 8192
rect 3434 8132 3438 8188
rect 3438 8132 3494 8188
rect 3494 8132 3498 8188
rect 3434 8128 3498 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 4929 8188 4993 8192
rect 4929 8132 4933 8188
rect 4933 8132 4989 8188
rect 4989 8132 4993 8188
rect 4929 8128 4993 8132
rect 6184 8188 6248 8192
rect 6184 8132 6188 8188
rect 6188 8132 6244 8188
rect 6244 8132 6248 8188
rect 6184 8128 6248 8132
rect 6264 8188 6328 8192
rect 6264 8132 6268 8188
rect 6268 8132 6324 8188
rect 6324 8132 6328 8188
rect 6264 8128 6328 8132
rect 6344 8188 6408 8192
rect 6344 8132 6348 8188
rect 6348 8132 6404 8188
rect 6404 8132 6408 8188
rect 6344 8128 6408 8132
rect 6424 8188 6488 8192
rect 6424 8132 6428 8188
rect 6428 8132 6484 8188
rect 6484 8132 6488 8188
rect 6424 8128 6488 8132
rect 2359 7644 2423 7648
rect 2359 7588 2363 7644
rect 2363 7588 2419 7644
rect 2419 7588 2423 7644
rect 2359 7584 2423 7588
rect 2439 7644 2503 7648
rect 2439 7588 2443 7644
rect 2443 7588 2499 7644
rect 2499 7588 2503 7644
rect 2439 7584 2503 7588
rect 2519 7644 2583 7648
rect 2519 7588 2523 7644
rect 2523 7588 2579 7644
rect 2579 7588 2583 7644
rect 2519 7584 2583 7588
rect 2599 7644 2663 7648
rect 2599 7588 2603 7644
rect 2603 7588 2659 7644
rect 2659 7588 2663 7644
rect 2599 7584 2663 7588
rect 3854 7644 3918 7648
rect 3854 7588 3858 7644
rect 3858 7588 3914 7644
rect 3914 7588 3918 7644
rect 3854 7584 3918 7588
rect 3934 7644 3998 7648
rect 3934 7588 3938 7644
rect 3938 7588 3994 7644
rect 3994 7588 3998 7644
rect 3934 7584 3998 7588
rect 4014 7644 4078 7648
rect 4014 7588 4018 7644
rect 4018 7588 4074 7644
rect 4074 7588 4078 7644
rect 4014 7584 4078 7588
rect 4094 7644 4158 7648
rect 4094 7588 4098 7644
rect 4098 7588 4154 7644
rect 4154 7588 4158 7644
rect 4094 7584 4158 7588
rect 5349 7644 5413 7648
rect 5349 7588 5353 7644
rect 5353 7588 5409 7644
rect 5409 7588 5413 7644
rect 5349 7584 5413 7588
rect 5429 7644 5493 7648
rect 5429 7588 5433 7644
rect 5433 7588 5489 7644
rect 5489 7588 5493 7644
rect 5429 7584 5493 7588
rect 5509 7644 5573 7648
rect 5509 7588 5513 7644
rect 5513 7588 5569 7644
rect 5569 7588 5573 7644
rect 5509 7584 5573 7588
rect 5589 7644 5653 7648
rect 5589 7588 5593 7644
rect 5593 7588 5649 7644
rect 5649 7588 5653 7644
rect 5589 7584 5653 7588
rect 6844 7644 6908 7648
rect 6844 7588 6848 7644
rect 6848 7588 6904 7644
rect 6904 7588 6908 7644
rect 6844 7584 6908 7588
rect 6924 7644 6988 7648
rect 6924 7588 6928 7644
rect 6928 7588 6984 7644
rect 6984 7588 6988 7644
rect 6924 7584 6988 7588
rect 7004 7644 7068 7648
rect 7004 7588 7008 7644
rect 7008 7588 7064 7644
rect 7064 7588 7068 7644
rect 7004 7584 7068 7588
rect 7084 7644 7148 7648
rect 7084 7588 7088 7644
rect 7088 7588 7144 7644
rect 7144 7588 7148 7644
rect 7084 7584 7148 7588
rect 1699 7100 1763 7104
rect 1699 7044 1703 7100
rect 1703 7044 1759 7100
rect 1759 7044 1763 7100
rect 1699 7040 1763 7044
rect 1779 7100 1843 7104
rect 1779 7044 1783 7100
rect 1783 7044 1839 7100
rect 1839 7044 1843 7100
rect 1779 7040 1843 7044
rect 1859 7100 1923 7104
rect 1859 7044 1863 7100
rect 1863 7044 1919 7100
rect 1919 7044 1923 7100
rect 1859 7040 1923 7044
rect 1939 7100 2003 7104
rect 1939 7044 1943 7100
rect 1943 7044 1999 7100
rect 1999 7044 2003 7100
rect 1939 7040 2003 7044
rect 3194 7100 3258 7104
rect 3194 7044 3198 7100
rect 3198 7044 3254 7100
rect 3254 7044 3258 7100
rect 3194 7040 3258 7044
rect 3274 7100 3338 7104
rect 3274 7044 3278 7100
rect 3278 7044 3334 7100
rect 3334 7044 3338 7100
rect 3274 7040 3338 7044
rect 3354 7100 3418 7104
rect 3354 7044 3358 7100
rect 3358 7044 3414 7100
rect 3414 7044 3418 7100
rect 3354 7040 3418 7044
rect 3434 7100 3498 7104
rect 3434 7044 3438 7100
rect 3438 7044 3494 7100
rect 3494 7044 3498 7100
rect 3434 7040 3498 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 4929 7100 4993 7104
rect 4929 7044 4933 7100
rect 4933 7044 4989 7100
rect 4989 7044 4993 7100
rect 4929 7040 4993 7044
rect 6184 7100 6248 7104
rect 6184 7044 6188 7100
rect 6188 7044 6244 7100
rect 6244 7044 6248 7100
rect 6184 7040 6248 7044
rect 6264 7100 6328 7104
rect 6264 7044 6268 7100
rect 6268 7044 6324 7100
rect 6324 7044 6328 7100
rect 6264 7040 6328 7044
rect 6344 7100 6408 7104
rect 6344 7044 6348 7100
rect 6348 7044 6404 7100
rect 6404 7044 6408 7100
rect 6344 7040 6408 7044
rect 6424 7100 6488 7104
rect 6424 7044 6428 7100
rect 6428 7044 6484 7100
rect 6484 7044 6488 7100
rect 6424 7040 6488 7044
rect 2359 6556 2423 6560
rect 2359 6500 2363 6556
rect 2363 6500 2419 6556
rect 2419 6500 2423 6556
rect 2359 6496 2423 6500
rect 2439 6556 2503 6560
rect 2439 6500 2443 6556
rect 2443 6500 2499 6556
rect 2499 6500 2503 6556
rect 2439 6496 2503 6500
rect 2519 6556 2583 6560
rect 2519 6500 2523 6556
rect 2523 6500 2579 6556
rect 2579 6500 2583 6556
rect 2519 6496 2583 6500
rect 2599 6556 2663 6560
rect 2599 6500 2603 6556
rect 2603 6500 2659 6556
rect 2659 6500 2663 6556
rect 2599 6496 2663 6500
rect 3854 6556 3918 6560
rect 3854 6500 3858 6556
rect 3858 6500 3914 6556
rect 3914 6500 3918 6556
rect 3854 6496 3918 6500
rect 3934 6556 3998 6560
rect 3934 6500 3938 6556
rect 3938 6500 3994 6556
rect 3994 6500 3998 6556
rect 3934 6496 3998 6500
rect 4014 6556 4078 6560
rect 4014 6500 4018 6556
rect 4018 6500 4074 6556
rect 4074 6500 4078 6556
rect 4014 6496 4078 6500
rect 4094 6556 4158 6560
rect 4094 6500 4098 6556
rect 4098 6500 4154 6556
rect 4154 6500 4158 6556
rect 4094 6496 4158 6500
rect 5349 6556 5413 6560
rect 5349 6500 5353 6556
rect 5353 6500 5409 6556
rect 5409 6500 5413 6556
rect 5349 6496 5413 6500
rect 5429 6556 5493 6560
rect 5429 6500 5433 6556
rect 5433 6500 5489 6556
rect 5489 6500 5493 6556
rect 5429 6496 5493 6500
rect 5509 6556 5573 6560
rect 5509 6500 5513 6556
rect 5513 6500 5569 6556
rect 5569 6500 5573 6556
rect 5509 6496 5573 6500
rect 5589 6556 5653 6560
rect 5589 6500 5593 6556
rect 5593 6500 5649 6556
rect 5649 6500 5653 6556
rect 5589 6496 5653 6500
rect 6844 6556 6908 6560
rect 6844 6500 6848 6556
rect 6848 6500 6904 6556
rect 6904 6500 6908 6556
rect 6844 6496 6908 6500
rect 6924 6556 6988 6560
rect 6924 6500 6928 6556
rect 6928 6500 6984 6556
rect 6984 6500 6988 6556
rect 6924 6496 6988 6500
rect 7004 6556 7068 6560
rect 7004 6500 7008 6556
rect 7008 6500 7064 6556
rect 7064 6500 7068 6556
rect 7004 6496 7068 6500
rect 7084 6556 7148 6560
rect 7084 6500 7088 6556
rect 7088 6500 7144 6556
rect 7144 6500 7148 6556
rect 7084 6496 7148 6500
rect 1699 6012 1763 6016
rect 1699 5956 1703 6012
rect 1703 5956 1759 6012
rect 1759 5956 1763 6012
rect 1699 5952 1763 5956
rect 1779 6012 1843 6016
rect 1779 5956 1783 6012
rect 1783 5956 1839 6012
rect 1839 5956 1843 6012
rect 1779 5952 1843 5956
rect 1859 6012 1923 6016
rect 1859 5956 1863 6012
rect 1863 5956 1919 6012
rect 1919 5956 1923 6012
rect 1859 5952 1923 5956
rect 1939 6012 2003 6016
rect 1939 5956 1943 6012
rect 1943 5956 1999 6012
rect 1999 5956 2003 6012
rect 1939 5952 2003 5956
rect 3194 6012 3258 6016
rect 3194 5956 3198 6012
rect 3198 5956 3254 6012
rect 3254 5956 3258 6012
rect 3194 5952 3258 5956
rect 3274 6012 3338 6016
rect 3274 5956 3278 6012
rect 3278 5956 3334 6012
rect 3334 5956 3338 6012
rect 3274 5952 3338 5956
rect 3354 6012 3418 6016
rect 3354 5956 3358 6012
rect 3358 5956 3414 6012
rect 3414 5956 3418 6012
rect 3354 5952 3418 5956
rect 3434 6012 3498 6016
rect 3434 5956 3438 6012
rect 3438 5956 3494 6012
rect 3494 5956 3498 6012
rect 3434 5952 3498 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 4929 6012 4993 6016
rect 4929 5956 4933 6012
rect 4933 5956 4989 6012
rect 4989 5956 4993 6012
rect 4929 5952 4993 5956
rect 6184 6012 6248 6016
rect 6184 5956 6188 6012
rect 6188 5956 6244 6012
rect 6244 5956 6248 6012
rect 6184 5952 6248 5956
rect 6264 6012 6328 6016
rect 6264 5956 6268 6012
rect 6268 5956 6324 6012
rect 6324 5956 6328 6012
rect 6264 5952 6328 5956
rect 6344 6012 6408 6016
rect 6344 5956 6348 6012
rect 6348 5956 6404 6012
rect 6404 5956 6408 6012
rect 6344 5952 6408 5956
rect 6424 6012 6488 6016
rect 6424 5956 6428 6012
rect 6428 5956 6484 6012
rect 6484 5956 6488 6012
rect 6424 5952 6488 5956
rect 2359 5468 2423 5472
rect 2359 5412 2363 5468
rect 2363 5412 2419 5468
rect 2419 5412 2423 5468
rect 2359 5408 2423 5412
rect 2439 5468 2503 5472
rect 2439 5412 2443 5468
rect 2443 5412 2499 5468
rect 2499 5412 2503 5468
rect 2439 5408 2503 5412
rect 2519 5468 2583 5472
rect 2519 5412 2523 5468
rect 2523 5412 2579 5468
rect 2579 5412 2583 5468
rect 2519 5408 2583 5412
rect 2599 5468 2663 5472
rect 2599 5412 2603 5468
rect 2603 5412 2659 5468
rect 2659 5412 2663 5468
rect 2599 5408 2663 5412
rect 3854 5468 3918 5472
rect 3854 5412 3858 5468
rect 3858 5412 3914 5468
rect 3914 5412 3918 5468
rect 3854 5408 3918 5412
rect 3934 5468 3998 5472
rect 3934 5412 3938 5468
rect 3938 5412 3994 5468
rect 3994 5412 3998 5468
rect 3934 5408 3998 5412
rect 4014 5468 4078 5472
rect 4014 5412 4018 5468
rect 4018 5412 4074 5468
rect 4074 5412 4078 5468
rect 4014 5408 4078 5412
rect 4094 5468 4158 5472
rect 4094 5412 4098 5468
rect 4098 5412 4154 5468
rect 4154 5412 4158 5468
rect 4094 5408 4158 5412
rect 5349 5468 5413 5472
rect 5349 5412 5353 5468
rect 5353 5412 5409 5468
rect 5409 5412 5413 5468
rect 5349 5408 5413 5412
rect 5429 5468 5493 5472
rect 5429 5412 5433 5468
rect 5433 5412 5489 5468
rect 5489 5412 5493 5468
rect 5429 5408 5493 5412
rect 5509 5468 5573 5472
rect 5509 5412 5513 5468
rect 5513 5412 5569 5468
rect 5569 5412 5573 5468
rect 5509 5408 5573 5412
rect 5589 5468 5653 5472
rect 5589 5412 5593 5468
rect 5593 5412 5649 5468
rect 5649 5412 5653 5468
rect 5589 5408 5653 5412
rect 6844 5468 6908 5472
rect 6844 5412 6848 5468
rect 6848 5412 6904 5468
rect 6904 5412 6908 5468
rect 6844 5408 6908 5412
rect 6924 5468 6988 5472
rect 6924 5412 6928 5468
rect 6928 5412 6984 5468
rect 6984 5412 6988 5468
rect 6924 5408 6988 5412
rect 7004 5468 7068 5472
rect 7004 5412 7008 5468
rect 7008 5412 7064 5468
rect 7064 5412 7068 5468
rect 7004 5408 7068 5412
rect 7084 5468 7148 5472
rect 7084 5412 7088 5468
rect 7088 5412 7144 5468
rect 7144 5412 7148 5468
rect 7084 5408 7148 5412
rect 1699 4924 1763 4928
rect 1699 4868 1703 4924
rect 1703 4868 1759 4924
rect 1759 4868 1763 4924
rect 1699 4864 1763 4868
rect 1779 4924 1843 4928
rect 1779 4868 1783 4924
rect 1783 4868 1839 4924
rect 1839 4868 1843 4924
rect 1779 4864 1843 4868
rect 1859 4924 1923 4928
rect 1859 4868 1863 4924
rect 1863 4868 1919 4924
rect 1919 4868 1923 4924
rect 1859 4864 1923 4868
rect 1939 4924 2003 4928
rect 1939 4868 1943 4924
rect 1943 4868 1999 4924
rect 1999 4868 2003 4924
rect 1939 4864 2003 4868
rect 3194 4924 3258 4928
rect 3194 4868 3198 4924
rect 3198 4868 3254 4924
rect 3254 4868 3258 4924
rect 3194 4864 3258 4868
rect 3274 4924 3338 4928
rect 3274 4868 3278 4924
rect 3278 4868 3334 4924
rect 3334 4868 3338 4924
rect 3274 4864 3338 4868
rect 3354 4924 3418 4928
rect 3354 4868 3358 4924
rect 3358 4868 3414 4924
rect 3414 4868 3418 4924
rect 3354 4864 3418 4868
rect 3434 4924 3498 4928
rect 3434 4868 3438 4924
rect 3438 4868 3494 4924
rect 3494 4868 3498 4924
rect 3434 4864 3498 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 4929 4924 4993 4928
rect 4929 4868 4933 4924
rect 4933 4868 4989 4924
rect 4989 4868 4993 4924
rect 4929 4864 4993 4868
rect 6184 4924 6248 4928
rect 6184 4868 6188 4924
rect 6188 4868 6244 4924
rect 6244 4868 6248 4924
rect 6184 4864 6248 4868
rect 6264 4924 6328 4928
rect 6264 4868 6268 4924
rect 6268 4868 6324 4924
rect 6324 4868 6328 4924
rect 6264 4864 6328 4868
rect 6344 4924 6408 4928
rect 6344 4868 6348 4924
rect 6348 4868 6404 4924
rect 6404 4868 6408 4924
rect 6344 4864 6408 4868
rect 6424 4924 6488 4928
rect 6424 4868 6428 4924
rect 6428 4868 6484 4924
rect 6484 4868 6488 4924
rect 6424 4864 6488 4868
rect 2359 4380 2423 4384
rect 2359 4324 2363 4380
rect 2363 4324 2419 4380
rect 2419 4324 2423 4380
rect 2359 4320 2423 4324
rect 2439 4380 2503 4384
rect 2439 4324 2443 4380
rect 2443 4324 2499 4380
rect 2499 4324 2503 4380
rect 2439 4320 2503 4324
rect 2519 4380 2583 4384
rect 2519 4324 2523 4380
rect 2523 4324 2579 4380
rect 2579 4324 2583 4380
rect 2519 4320 2583 4324
rect 2599 4380 2663 4384
rect 2599 4324 2603 4380
rect 2603 4324 2659 4380
rect 2659 4324 2663 4380
rect 2599 4320 2663 4324
rect 3854 4380 3918 4384
rect 3854 4324 3858 4380
rect 3858 4324 3914 4380
rect 3914 4324 3918 4380
rect 3854 4320 3918 4324
rect 3934 4380 3998 4384
rect 3934 4324 3938 4380
rect 3938 4324 3994 4380
rect 3994 4324 3998 4380
rect 3934 4320 3998 4324
rect 4014 4380 4078 4384
rect 4014 4324 4018 4380
rect 4018 4324 4074 4380
rect 4074 4324 4078 4380
rect 4014 4320 4078 4324
rect 4094 4380 4158 4384
rect 4094 4324 4098 4380
rect 4098 4324 4154 4380
rect 4154 4324 4158 4380
rect 4094 4320 4158 4324
rect 5349 4380 5413 4384
rect 5349 4324 5353 4380
rect 5353 4324 5409 4380
rect 5409 4324 5413 4380
rect 5349 4320 5413 4324
rect 5429 4380 5493 4384
rect 5429 4324 5433 4380
rect 5433 4324 5489 4380
rect 5489 4324 5493 4380
rect 5429 4320 5493 4324
rect 5509 4380 5573 4384
rect 5509 4324 5513 4380
rect 5513 4324 5569 4380
rect 5569 4324 5573 4380
rect 5509 4320 5573 4324
rect 5589 4380 5653 4384
rect 5589 4324 5593 4380
rect 5593 4324 5649 4380
rect 5649 4324 5653 4380
rect 5589 4320 5653 4324
rect 6844 4380 6908 4384
rect 6844 4324 6848 4380
rect 6848 4324 6904 4380
rect 6904 4324 6908 4380
rect 6844 4320 6908 4324
rect 6924 4380 6988 4384
rect 6924 4324 6928 4380
rect 6928 4324 6984 4380
rect 6984 4324 6988 4380
rect 6924 4320 6988 4324
rect 7004 4380 7068 4384
rect 7004 4324 7008 4380
rect 7008 4324 7064 4380
rect 7064 4324 7068 4380
rect 7004 4320 7068 4324
rect 7084 4380 7148 4384
rect 7084 4324 7088 4380
rect 7088 4324 7144 4380
rect 7144 4324 7148 4380
rect 7084 4320 7148 4324
rect 1699 3836 1763 3840
rect 1699 3780 1703 3836
rect 1703 3780 1759 3836
rect 1759 3780 1763 3836
rect 1699 3776 1763 3780
rect 1779 3836 1843 3840
rect 1779 3780 1783 3836
rect 1783 3780 1839 3836
rect 1839 3780 1843 3836
rect 1779 3776 1843 3780
rect 1859 3836 1923 3840
rect 1859 3780 1863 3836
rect 1863 3780 1919 3836
rect 1919 3780 1923 3836
rect 1859 3776 1923 3780
rect 1939 3836 2003 3840
rect 1939 3780 1943 3836
rect 1943 3780 1999 3836
rect 1999 3780 2003 3836
rect 1939 3776 2003 3780
rect 3194 3836 3258 3840
rect 3194 3780 3198 3836
rect 3198 3780 3254 3836
rect 3254 3780 3258 3836
rect 3194 3776 3258 3780
rect 3274 3836 3338 3840
rect 3274 3780 3278 3836
rect 3278 3780 3334 3836
rect 3334 3780 3338 3836
rect 3274 3776 3338 3780
rect 3354 3836 3418 3840
rect 3354 3780 3358 3836
rect 3358 3780 3414 3836
rect 3414 3780 3418 3836
rect 3354 3776 3418 3780
rect 3434 3836 3498 3840
rect 3434 3780 3438 3836
rect 3438 3780 3494 3836
rect 3494 3780 3498 3836
rect 3434 3776 3498 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 4929 3836 4993 3840
rect 4929 3780 4933 3836
rect 4933 3780 4989 3836
rect 4989 3780 4993 3836
rect 4929 3776 4993 3780
rect 6184 3836 6248 3840
rect 6184 3780 6188 3836
rect 6188 3780 6244 3836
rect 6244 3780 6248 3836
rect 6184 3776 6248 3780
rect 6264 3836 6328 3840
rect 6264 3780 6268 3836
rect 6268 3780 6324 3836
rect 6324 3780 6328 3836
rect 6264 3776 6328 3780
rect 6344 3836 6408 3840
rect 6344 3780 6348 3836
rect 6348 3780 6404 3836
rect 6404 3780 6408 3836
rect 6344 3776 6408 3780
rect 6424 3836 6488 3840
rect 6424 3780 6428 3836
rect 6428 3780 6484 3836
rect 6484 3780 6488 3836
rect 6424 3776 6488 3780
rect 2359 3292 2423 3296
rect 2359 3236 2363 3292
rect 2363 3236 2419 3292
rect 2419 3236 2423 3292
rect 2359 3232 2423 3236
rect 2439 3292 2503 3296
rect 2439 3236 2443 3292
rect 2443 3236 2499 3292
rect 2499 3236 2503 3292
rect 2439 3232 2503 3236
rect 2519 3292 2583 3296
rect 2519 3236 2523 3292
rect 2523 3236 2579 3292
rect 2579 3236 2583 3292
rect 2519 3232 2583 3236
rect 2599 3292 2663 3296
rect 2599 3236 2603 3292
rect 2603 3236 2659 3292
rect 2659 3236 2663 3292
rect 2599 3232 2663 3236
rect 3854 3292 3918 3296
rect 3854 3236 3858 3292
rect 3858 3236 3914 3292
rect 3914 3236 3918 3292
rect 3854 3232 3918 3236
rect 3934 3292 3998 3296
rect 3934 3236 3938 3292
rect 3938 3236 3994 3292
rect 3994 3236 3998 3292
rect 3934 3232 3998 3236
rect 4014 3292 4078 3296
rect 4014 3236 4018 3292
rect 4018 3236 4074 3292
rect 4074 3236 4078 3292
rect 4014 3232 4078 3236
rect 4094 3292 4158 3296
rect 4094 3236 4098 3292
rect 4098 3236 4154 3292
rect 4154 3236 4158 3292
rect 4094 3232 4158 3236
rect 5349 3292 5413 3296
rect 5349 3236 5353 3292
rect 5353 3236 5409 3292
rect 5409 3236 5413 3292
rect 5349 3232 5413 3236
rect 5429 3292 5493 3296
rect 5429 3236 5433 3292
rect 5433 3236 5489 3292
rect 5489 3236 5493 3292
rect 5429 3232 5493 3236
rect 5509 3292 5573 3296
rect 5509 3236 5513 3292
rect 5513 3236 5569 3292
rect 5569 3236 5573 3292
rect 5509 3232 5573 3236
rect 5589 3292 5653 3296
rect 5589 3236 5593 3292
rect 5593 3236 5649 3292
rect 5649 3236 5653 3292
rect 5589 3232 5653 3236
rect 6844 3292 6908 3296
rect 6844 3236 6848 3292
rect 6848 3236 6904 3292
rect 6904 3236 6908 3292
rect 6844 3232 6908 3236
rect 6924 3292 6988 3296
rect 6924 3236 6928 3292
rect 6928 3236 6984 3292
rect 6984 3236 6988 3292
rect 6924 3232 6988 3236
rect 7004 3292 7068 3296
rect 7004 3236 7008 3292
rect 7008 3236 7064 3292
rect 7064 3236 7068 3292
rect 7004 3232 7068 3236
rect 7084 3292 7148 3296
rect 7084 3236 7088 3292
rect 7088 3236 7144 3292
rect 7144 3236 7148 3292
rect 7084 3232 7148 3236
rect 1699 2748 1763 2752
rect 1699 2692 1703 2748
rect 1703 2692 1759 2748
rect 1759 2692 1763 2748
rect 1699 2688 1763 2692
rect 1779 2748 1843 2752
rect 1779 2692 1783 2748
rect 1783 2692 1839 2748
rect 1839 2692 1843 2748
rect 1779 2688 1843 2692
rect 1859 2748 1923 2752
rect 1859 2692 1863 2748
rect 1863 2692 1919 2748
rect 1919 2692 1923 2748
rect 1859 2688 1923 2692
rect 1939 2748 2003 2752
rect 1939 2692 1943 2748
rect 1943 2692 1999 2748
rect 1999 2692 2003 2748
rect 1939 2688 2003 2692
rect 3194 2748 3258 2752
rect 3194 2692 3198 2748
rect 3198 2692 3254 2748
rect 3254 2692 3258 2748
rect 3194 2688 3258 2692
rect 3274 2748 3338 2752
rect 3274 2692 3278 2748
rect 3278 2692 3334 2748
rect 3334 2692 3338 2748
rect 3274 2688 3338 2692
rect 3354 2748 3418 2752
rect 3354 2692 3358 2748
rect 3358 2692 3414 2748
rect 3414 2692 3418 2748
rect 3354 2688 3418 2692
rect 3434 2748 3498 2752
rect 3434 2692 3438 2748
rect 3438 2692 3494 2748
rect 3494 2692 3498 2748
rect 3434 2688 3498 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 4929 2748 4993 2752
rect 4929 2692 4933 2748
rect 4933 2692 4989 2748
rect 4989 2692 4993 2748
rect 4929 2688 4993 2692
rect 6184 2748 6248 2752
rect 6184 2692 6188 2748
rect 6188 2692 6244 2748
rect 6244 2692 6248 2748
rect 6184 2688 6248 2692
rect 6264 2748 6328 2752
rect 6264 2692 6268 2748
rect 6268 2692 6324 2748
rect 6324 2692 6328 2748
rect 6264 2688 6328 2692
rect 6344 2748 6408 2752
rect 6344 2692 6348 2748
rect 6348 2692 6404 2748
rect 6404 2692 6408 2748
rect 6344 2688 6408 2692
rect 6424 2748 6488 2752
rect 6424 2692 6428 2748
rect 6428 2692 6484 2748
rect 6484 2692 6488 2748
rect 6424 2688 6488 2692
rect 2359 2204 2423 2208
rect 2359 2148 2363 2204
rect 2363 2148 2419 2204
rect 2419 2148 2423 2204
rect 2359 2144 2423 2148
rect 2439 2204 2503 2208
rect 2439 2148 2443 2204
rect 2443 2148 2499 2204
rect 2499 2148 2503 2204
rect 2439 2144 2503 2148
rect 2519 2204 2583 2208
rect 2519 2148 2523 2204
rect 2523 2148 2579 2204
rect 2579 2148 2583 2204
rect 2519 2144 2583 2148
rect 2599 2204 2663 2208
rect 2599 2148 2603 2204
rect 2603 2148 2659 2204
rect 2659 2148 2663 2204
rect 2599 2144 2663 2148
rect 3854 2204 3918 2208
rect 3854 2148 3858 2204
rect 3858 2148 3914 2204
rect 3914 2148 3918 2204
rect 3854 2144 3918 2148
rect 3934 2204 3998 2208
rect 3934 2148 3938 2204
rect 3938 2148 3994 2204
rect 3994 2148 3998 2204
rect 3934 2144 3998 2148
rect 4014 2204 4078 2208
rect 4014 2148 4018 2204
rect 4018 2148 4074 2204
rect 4074 2148 4078 2204
rect 4014 2144 4078 2148
rect 4094 2204 4158 2208
rect 4094 2148 4098 2204
rect 4098 2148 4154 2204
rect 4154 2148 4158 2204
rect 4094 2144 4158 2148
rect 5349 2204 5413 2208
rect 5349 2148 5353 2204
rect 5353 2148 5409 2204
rect 5409 2148 5413 2204
rect 5349 2144 5413 2148
rect 5429 2204 5493 2208
rect 5429 2148 5433 2204
rect 5433 2148 5489 2204
rect 5489 2148 5493 2204
rect 5429 2144 5493 2148
rect 5509 2204 5573 2208
rect 5509 2148 5513 2204
rect 5513 2148 5569 2204
rect 5569 2148 5573 2204
rect 5509 2144 5573 2148
rect 5589 2204 5653 2208
rect 5589 2148 5593 2204
rect 5593 2148 5649 2204
rect 5649 2148 5653 2204
rect 5589 2144 5653 2148
rect 6844 2204 6908 2208
rect 6844 2148 6848 2204
rect 6848 2148 6904 2204
rect 6904 2148 6908 2204
rect 6844 2144 6908 2148
rect 6924 2204 6988 2208
rect 6924 2148 6928 2204
rect 6928 2148 6984 2204
rect 6984 2148 6988 2204
rect 6924 2144 6988 2148
rect 7004 2204 7068 2208
rect 7004 2148 7008 2204
rect 7008 2148 7064 2204
rect 7064 2148 7068 2204
rect 7004 2144 7068 2148
rect 7084 2204 7148 2208
rect 7084 2148 7088 2204
rect 7088 2148 7144 2204
rect 7144 2148 7148 2204
rect 7084 2144 7148 2148
<< metal4 >>
rect 1691 8192 2011 8208
rect 1691 8128 1699 8192
rect 1763 8128 1779 8192
rect 1843 8128 1859 8192
rect 1923 8128 1939 8192
rect 2003 8128 2011 8192
rect 1691 7526 2011 8128
rect 1691 7290 1733 7526
rect 1969 7290 2011 7526
rect 1691 7104 2011 7290
rect 1691 7040 1699 7104
rect 1763 7040 1779 7104
rect 1843 7040 1859 7104
rect 1923 7040 1939 7104
rect 2003 7040 2011 7104
rect 1691 6031 2011 7040
rect 1691 6016 1733 6031
rect 1969 6016 2011 6031
rect 1691 5952 1699 6016
rect 2003 5952 2011 6016
rect 1691 5795 1733 5952
rect 1969 5795 2011 5952
rect 1691 4928 2011 5795
rect 1691 4864 1699 4928
rect 1763 4864 1779 4928
rect 1843 4864 1859 4928
rect 1923 4864 1939 4928
rect 2003 4864 2011 4928
rect 1691 4536 2011 4864
rect 1691 4300 1733 4536
rect 1969 4300 2011 4536
rect 1691 3840 2011 4300
rect 1691 3776 1699 3840
rect 1763 3776 1779 3840
rect 1843 3776 1859 3840
rect 1923 3776 1939 3840
rect 2003 3776 2011 3840
rect 1691 3041 2011 3776
rect 1691 2805 1733 3041
rect 1969 2805 2011 3041
rect 1691 2752 2011 2805
rect 1691 2688 1699 2752
rect 1763 2688 1779 2752
rect 1843 2688 1859 2752
rect 1923 2688 1939 2752
rect 2003 2688 2011 2752
rect 1691 2128 2011 2688
rect 2351 8186 2671 8228
rect 2351 7950 2393 8186
rect 2629 7950 2671 8186
rect 2351 7648 2671 7950
rect 2351 7584 2359 7648
rect 2423 7584 2439 7648
rect 2503 7584 2519 7648
rect 2583 7584 2599 7648
rect 2663 7584 2671 7648
rect 2351 6691 2671 7584
rect 2351 6560 2393 6691
rect 2629 6560 2671 6691
rect 2351 6496 2359 6560
rect 2663 6496 2671 6560
rect 2351 6455 2393 6496
rect 2629 6455 2671 6496
rect 2351 5472 2671 6455
rect 2351 5408 2359 5472
rect 2423 5408 2439 5472
rect 2503 5408 2519 5472
rect 2583 5408 2599 5472
rect 2663 5408 2671 5472
rect 2351 5196 2671 5408
rect 2351 4960 2393 5196
rect 2629 4960 2671 5196
rect 2351 4384 2671 4960
rect 2351 4320 2359 4384
rect 2423 4320 2439 4384
rect 2503 4320 2519 4384
rect 2583 4320 2599 4384
rect 2663 4320 2671 4384
rect 2351 3701 2671 4320
rect 2351 3465 2393 3701
rect 2629 3465 2671 3701
rect 2351 3296 2671 3465
rect 2351 3232 2359 3296
rect 2423 3232 2439 3296
rect 2503 3232 2519 3296
rect 2583 3232 2599 3296
rect 2663 3232 2671 3296
rect 2351 2208 2671 3232
rect 2351 2144 2359 2208
rect 2423 2144 2439 2208
rect 2503 2144 2519 2208
rect 2583 2144 2599 2208
rect 2663 2144 2671 2208
rect 2351 2128 2671 2144
rect 3186 8192 3506 8208
rect 3186 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3434 8192
rect 3498 8128 3506 8192
rect 3186 7526 3506 8128
rect 3186 7290 3228 7526
rect 3464 7290 3506 7526
rect 3186 7104 3506 7290
rect 3186 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3434 7104
rect 3498 7040 3506 7104
rect 3186 6031 3506 7040
rect 3186 6016 3228 6031
rect 3464 6016 3506 6031
rect 3186 5952 3194 6016
rect 3498 5952 3506 6016
rect 3186 5795 3228 5952
rect 3464 5795 3506 5952
rect 3186 4928 3506 5795
rect 3186 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3434 4928
rect 3498 4864 3506 4928
rect 3186 4536 3506 4864
rect 3186 4300 3228 4536
rect 3464 4300 3506 4536
rect 3186 3840 3506 4300
rect 3186 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3434 3840
rect 3498 3776 3506 3840
rect 3186 3041 3506 3776
rect 3186 2805 3228 3041
rect 3464 2805 3506 3041
rect 3186 2752 3506 2805
rect 3186 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3434 2752
rect 3498 2688 3506 2752
rect 3186 2128 3506 2688
rect 3846 8186 4166 8228
rect 3846 7950 3888 8186
rect 4124 7950 4166 8186
rect 3846 7648 4166 7950
rect 3846 7584 3854 7648
rect 3918 7584 3934 7648
rect 3998 7584 4014 7648
rect 4078 7584 4094 7648
rect 4158 7584 4166 7648
rect 3846 6691 4166 7584
rect 3846 6560 3888 6691
rect 4124 6560 4166 6691
rect 3846 6496 3854 6560
rect 4158 6496 4166 6560
rect 3846 6455 3888 6496
rect 4124 6455 4166 6496
rect 3846 5472 4166 6455
rect 3846 5408 3854 5472
rect 3918 5408 3934 5472
rect 3998 5408 4014 5472
rect 4078 5408 4094 5472
rect 4158 5408 4166 5472
rect 3846 5196 4166 5408
rect 3846 4960 3888 5196
rect 4124 4960 4166 5196
rect 3846 4384 4166 4960
rect 3846 4320 3854 4384
rect 3918 4320 3934 4384
rect 3998 4320 4014 4384
rect 4078 4320 4094 4384
rect 4158 4320 4166 4384
rect 3846 3701 4166 4320
rect 3846 3465 3888 3701
rect 4124 3465 4166 3701
rect 3846 3296 4166 3465
rect 3846 3232 3854 3296
rect 3918 3232 3934 3296
rect 3998 3232 4014 3296
rect 4078 3232 4094 3296
rect 4158 3232 4166 3296
rect 3846 2208 4166 3232
rect 3846 2144 3854 2208
rect 3918 2144 3934 2208
rect 3998 2144 4014 2208
rect 4078 2144 4094 2208
rect 4158 2144 4166 2208
rect 3846 2128 4166 2144
rect 4681 8192 5001 8208
rect 4681 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4929 8192
rect 4993 8128 5001 8192
rect 4681 7526 5001 8128
rect 4681 7290 4723 7526
rect 4959 7290 5001 7526
rect 4681 7104 5001 7290
rect 4681 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4929 7104
rect 4993 7040 5001 7104
rect 4681 6031 5001 7040
rect 4681 6016 4723 6031
rect 4959 6016 5001 6031
rect 4681 5952 4689 6016
rect 4993 5952 5001 6016
rect 4681 5795 4723 5952
rect 4959 5795 5001 5952
rect 4681 4928 5001 5795
rect 4681 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4929 4928
rect 4993 4864 5001 4928
rect 4681 4536 5001 4864
rect 4681 4300 4723 4536
rect 4959 4300 5001 4536
rect 4681 3840 5001 4300
rect 4681 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4929 3840
rect 4993 3776 5001 3840
rect 4681 3041 5001 3776
rect 4681 2805 4723 3041
rect 4959 2805 5001 3041
rect 4681 2752 5001 2805
rect 4681 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4929 2752
rect 4993 2688 5001 2752
rect 4681 2128 5001 2688
rect 5341 8186 5661 8228
rect 5341 7950 5383 8186
rect 5619 7950 5661 8186
rect 5341 7648 5661 7950
rect 5341 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5589 7648
rect 5653 7584 5661 7648
rect 5341 6691 5661 7584
rect 5341 6560 5383 6691
rect 5619 6560 5661 6691
rect 5341 6496 5349 6560
rect 5653 6496 5661 6560
rect 5341 6455 5383 6496
rect 5619 6455 5661 6496
rect 5341 5472 5661 6455
rect 5341 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5589 5472
rect 5653 5408 5661 5472
rect 5341 5196 5661 5408
rect 5341 4960 5383 5196
rect 5619 4960 5661 5196
rect 5341 4384 5661 4960
rect 5341 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5589 4384
rect 5653 4320 5661 4384
rect 5341 3701 5661 4320
rect 5341 3465 5383 3701
rect 5619 3465 5661 3701
rect 5341 3296 5661 3465
rect 5341 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5589 3296
rect 5653 3232 5661 3296
rect 5341 2208 5661 3232
rect 5341 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5589 2208
rect 5653 2144 5661 2208
rect 5341 2128 5661 2144
rect 6176 8192 6496 8208
rect 6176 8128 6184 8192
rect 6248 8128 6264 8192
rect 6328 8128 6344 8192
rect 6408 8128 6424 8192
rect 6488 8128 6496 8192
rect 6176 7526 6496 8128
rect 6176 7290 6218 7526
rect 6454 7290 6496 7526
rect 6176 7104 6496 7290
rect 6176 7040 6184 7104
rect 6248 7040 6264 7104
rect 6328 7040 6344 7104
rect 6408 7040 6424 7104
rect 6488 7040 6496 7104
rect 6176 6031 6496 7040
rect 6176 6016 6218 6031
rect 6454 6016 6496 6031
rect 6176 5952 6184 6016
rect 6488 5952 6496 6016
rect 6176 5795 6218 5952
rect 6454 5795 6496 5952
rect 6176 4928 6496 5795
rect 6176 4864 6184 4928
rect 6248 4864 6264 4928
rect 6328 4864 6344 4928
rect 6408 4864 6424 4928
rect 6488 4864 6496 4928
rect 6176 4536 6496 4864
rect 6176 4300 6218 4536
rect 6454 4300 6496 4536
rect 6176 3840 6496 4300
rect 6176 3776 6184 3840
rect 6248 3776 6264 3840
rect 6328 3776 6344 3840
rect 6408 3776 6424 3840
rect 6488 3776 6496 3840
rect 6176 3041 6496 3776
rect 6176 2805 6218 3041
rect 6454 2805 6496 3041
rect 6176 2752 6496 2805
rect 6176 2688 6184 2752
rect 6248 2688 6264 2752
rect 6328 2688 6344 2752
rect 6408 2688 6424 2752
rect 6488 2688 6496 2752
rect 6176 2128 6496 2688
rect 6836 8186 7156 8228
rect 6836 7950 6878 8186
rect 7114 7950 7156 8186
rect 6836 7648 7156 7950
rect 6836 7584 6844 7648
rect 6908 7584 6924 7648
rect 6988 7584 7004 7648
rect 7068 7584 7084 7648
rect 7148 7584 7156 7648
rect 6836 6691 7156 7584
rect 6836 6560 6878 6691
rect 7114 6560 7156 6691
rect 6836 6496 6844 6560
rect 7148 6496 7156 6560
rect 6836 6455 6878 6496
rect 7114 6455 7156 6496
rect 6836 5472 7156 6455
rect 6836 5408 6844 5472
rect 6908 5408 6924 5472
rect 6988 5408 7004 5472
rect 7068 5408 7084 5472
rect 7148 5408 7156 5472
rect 6836 5196 7156 5408
rect 6836 4960 6878 5196
rect 7114 4960 7156 5196
rect 6836 4384 7156 4960
rect 6836 4320 6844 4384
rect 6908 4320 6924 4384
rect 6988 4320 7004 4384
rect 7068 4320 7084 4384
rect 7148 4320 7156 4384
rect 6836 3701 7156 4320
rect 6836 3465 6878 3701
rect 7114 3465 7156 3701
rect 6836 3296 7156 3465
rect 6836 3232 6844 3296
rect 6908 3232 6924 3296
rect 6988 3232 7004 3296
rect 7068 3232 7084 3296
rect 7148 3232 7156 3296
rect 6836 2208 7156 3232
rect 6836 2144 6844 2208
rect 6908 2144 6924 2208
rect 6988 2144 7004 2208
rect 7068 2144 7084 2208
rect 7148 2144 7156 2208
rect 6836 2128 7156 2144
<< via4 >>
rect 1733 7290 1969 7526
rect 1733 6016 1969 6031
rect 1733 5952 1763 6016
rect 1763 5952 1779 6016
rect 1779 5952 1843 6016
rect 1843 5952 1859 6016
rect 1859 5952 1923 6016
rect 1923 5952 1939 6016
rect 1939 5952 1969 6016
rect 1733 5795 1969 5952
rect 1733 4300 1969 4536
rect 1733 2805 1969 3041
rect 2393 7950 2629 8186
rect 2393 6560 2629 6691
rect 2393 6496 2423 6560
rect 2423 6496 2439 6560
rect 2439 6496 2503 6560
rect 2503 6496 2519 6560
rect 2519 6496 2583 6560
rect 2583 6496 2599 6560
rect 2599 6496 2629 6560
rect 2393 6455 2629 6496
rect 2393 4960 2629 5196
rect 2393 3465 2629 3701
rect 3228 7290 3464 7526
rect 3228 6016 3464 6031
rect 3228 5952 3258 6016
rect 3258 5952 3274 6016
rect 3274 5952 3338 6016
rect 3338 5952 3354 6016
rect 3354 5952 3418 6016
rect 3418 5952 3434 6016
rect 3434 5952 3464 6016
rect 3228 5795 3464 5952
rect 3228 4300 3464 4536
rect 3228 2805 3464 3041
rect 3888 7950 4124 8186
rect 3888 6560 4124 6691
rect 3888 6496 3918 6560
rect 3918 6496 3934 6560
rect 3934 6496 3998 6560
rect 3998 6496 4014 6560
rect 4014 6496 4078 6560
rect 4078 6496 4094 6560
rect 4094 6496 4124 6560
rect 3888 6455 4124 6496
rect 3888 4960 4124 5196
rect 3888 3465 4124 3701
rect 4723 7290 4959 7526
rect 4723 6016 4959 6031
rect 4723 5952 4753 6016
rect 4753 5952 4769 6016
rect 4769 5952 4833 6016
rect 4833 5952 4849 6016
rect 4849 5952 4913 6016
rect 4913 5952 4929 6016
rect 4929 5952 4959 6016
rect 4723 5795 4959 5952
rect 4723 4300 4959 4536
rect 4723 2805 4959 3041
rect 5383 7950 5619 8186
rect 5383 6560 5619 6691
rect 5383 6496 5413 6560
rect 5413 6496 5429 6560
rect 5429 6496 5493 6560
rect 5493 6496 5509 6560
rect 5509 6496 5573 6560
rect 5573 6496 5589 6560
rect 5589 6496 5619 6560
rect 5383 6455 5619 6496
rect 5383 4960 5619 5196
rect 5383 3465 5619 3701
rect 6218 7290 6454 7526
rect 6218 6016 6454 6031
rect 6218 5952 6248 6016
rect 6248 5952 6264 6016
rect 6264 5952 6328 6016
rect 6328 5952 6344 6016
rect 6344 5952 6408 6016
rect 6408 5952 6424 6016
rect 6424 5952 6454 6016
rect 6218 5795 6454 5952
rect 6218 4300 6454 4536
rect 6218 2805 6454 3041
rect 6878 7950 7114 8186
rect 6878 6560 7114 6691
rect 6878 6496 6908 6560
rect 6908 6496 6924 6560
rect 6924 6496 6988 6560
rect 6988 6496 7004 6560
rect 7004 6496 7068 6560
rect 7068 6496 7084 6560
rect 7084 6496 7114 6560
rect 6878 6455 7114 6496
rect 6878 4960 7114 5196
rect 6878 3465 7114 3701
<< metal5 >>
rect 1056 8186 7156 8228
rect 1056 7950 2393 8186
rect 2629 7950 3888 8186
rect 4124 7950 5383 8186
rect 5619 7950 6878 8186
rect 7114 7950 7156 8186
rect 1056 7908 7156 7950
rect 1056 7526 7132 7568
rect 1056 7290 1733 7526
rect 1969 7290 3228 7526
rect 3464 7290 4723 7526
rect 4959 7290 6218 7526
rect 6454 7290 7132 7526
rect 1056 7248 7132 7290
rect 1056 6691 7156 6733
rect 1056 6455 2393 6691
rect 2629 6455 3888 6691
rect 4124 6455 5383 6691
rect 5619 6455 6878 6691
rect 7114 6455 7156 6691
rect 1056 6413 7156 6455
rect 1056 6031 7132 6073
rect 1056 5795 1733 6031
rect 1969 5795 3228 6031
rect 3464 5795 4723 6031
rect 4959 5795 6218 6031
rect 6454 5795 7132 6031
rect 1056 5753 7132 5795
rect 1056 5196 7156 5238
rect 1056 4960 2393 5196
rect 2629 4960 3888 5196
rect 4124 4960 5383 5196
rect 5619 4960 6878 5196
rect 7114 4960 7156 5196
rect 1056 4918 7156 4960
rect 1056 4536 7132 4578
rect 1056 4300 1733 4536
rect 1969 4300 3228 4536
rect 3464 4300 4723 4536
rect 4959 4300 6218 4536
rect 6454 4300 7132 4536
rect 1056 4258 7132 4300
rect 1056 3701 7156 3743
rect 1056 3465 2393 3701
rect 2629 3465 3888 3701
rect 4124 3465 5383 3701
rect 5619 3465 6878 3701
rect 7114 3465 7156 3701
rect 1056 3423 7156 3465
rect 1056 3041 7132 3083
rect 1056 2805 1733 3041
rect 1969 2805 3228 3041
rect 3464 2805 4723 3041
rect 4959 2805 6218 3041
rect 6454 2805 7132 3041
rect 1056 2763 7132 2805
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_12
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1676037725
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1676037725
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1676037725
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1676037725
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_13
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1676037725
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1676037725
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1676037725
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1676037725
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1676037725
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1676037725
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6072 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1676037725
transform 1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1676037725
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 1676037725
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1676037725
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1676037725
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1676037725
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1676037725
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1676037725
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1676037725
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1676037725
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1676037725
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1676037725
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_45
timestamp 1676037725
transform 1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1676037725
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1676037725
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_60
timestamp 1676037725
transform 1 0 6624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1676037725
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1676037725
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1676037725
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_34
timestamp 1676037725
transform 1 0 4232 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1676037725
transform 1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_54
timestamp 1676037725
transform 1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1676037725
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1676037725
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5704 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4508 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _29_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _31_
timestamp 1676037725
transform 1 0 4784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1676037725
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _33_
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _34_
timestamp 1676037725
transform 1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1676037725
transform -1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _36_
timestamp 1676037725
transform -1 0 5336 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _37_
timestamp 1676037725
transform 1 0 4876 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1676037725
transform -1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _39_
timestamp 1676037725
transform 1 0 1656 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _40__1
timestamp 1676037725
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _41_
timestamp 1676037725
transform -1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _42_
timestamp 1676037725
transform 1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _43_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _44_
timestamp 1676037725
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _45_
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _46__2
timestamp 1676037725
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _47_
timestamp 1676037725
transform -1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _48_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _49_
timestamp 1676037725
transform 1 0 5152 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _50_
timestamp 1676037725
transform -1 0 6072 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _51_
timestamp 1676037725
transform 1 0 3312 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _52_
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _53_
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _54_
timestamp 1676037725
transform -1 0 3496 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _55_
timestamp 1676037725
transform -1 0 3496 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 3404 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform 1 0 2576 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform -1 0 4232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1676037725
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1676037725
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1676037725
transform -1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1676037725
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1676037725
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1676037725
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
<< labels >>
flabel metal4 s 2351 2128 2671 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3846 2128 4166 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5341 2128 5661 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6836 2128 7156 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3423 7156 3743 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4918 7156 5238 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6413 7156 6733 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7908 7156 8228 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1691 2128 2011 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3186 2128 3506 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4681 2128 5001 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6176 2128 6496 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2763 7132 3083 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4258 7132 4578 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5753 7132 6073 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7248 7132 7568 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 7458 1368 8258 1488 0 FreeSans 480 0 0 0 q[0]
port 3 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 q[1]
port 4 nsew signal tristate
flabel metal2 s 6458 9602 6514 10402 0 FreeSans 224 90 0 0 q[2]
port 5 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 q[3]
port 6 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 qb[0]
port 7 nsew signal tristate
flabel metal3 s 7458 8848 8258 8968 0 FreeSans 480 0 0 0 qb[1]
port 8 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 qb[2]
port 9 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 qb[3]
port 10 nsew signal tristate
flabel metal2 s 3238 9602 3294 10402 0 FreeSans 224 90 0 0 rst
port 11 nsew signal input
flabel metal3 s 7458 5448 8258 5568 0 FreeSans 480 0 0 0 t
port 12 nsew signal input
rlabel via1 4130 7616 4130 7616 0 VGND
rlabel metal1 4094 8160 4094 8160 0 VPWR
rlabel metal2 4186 3740 4186 3740 0 _01_
rlabel metal1 5980 4794 5980 4794 0 _02_
rlabel metal1 3128 2958 3128 2958 0 _03_
rlabel metal2 2070 3604 2070 3604 0 _04_
rlabel metal1 2990 2618 2990 2618 0 _05_
rlabel metal1 3450 6324 3450 6324 0 _07_
rlabel metal1 1978 3706 1978 3706 0 _08_
rlabel metal1 5336 3162 5336 3162 0 _09_
rlabel metal2 5290 6086 5290 6086 0 _10_
rlabel metal2 3082 4046 3082 4046 0 _11_
rlabel metal1 3818 2618 3818 2618 0 _12_
rlabel via1 4273 4590 4273 4590 0 _13_
rlabel metal2 5842 4352 5842 4352 0 _14_
rlabel metal2 2898 5542 2898 5542 0 _15_
rlabel metal1 2024 4590 2024 4590 0 _16_
rlabel metal2 2254 3553 2254 3553 0 _17_
rlabel metal2 1978 3162 1978 3162 0 _18_
rlabel metal1 5244 5338 5244 5338 0 _19_
rlabel metal2 6026 3196 6026 3196 0 _20_
rlabel metal1 4738 5338 4738 5338 0 _21_
rlabel metal2 2714 4454 2714 4454 0 _22_
rlabel metal2 5198 3468 5198 3468 0 _23_
rlabel metal3 820 6868 820 6868 0 clk
rlabel metal1 3220 7786 3220 7786 0 clknet_0_clk
rlabel metal1 2208 7378 2208 7378 0 clknet_1_0__leaf_clk
rlabel metal1 3818 6290 3818 6290 0 clknet_1_1__leaf_clk
rlabel metal2 4462 7242 4462 7242 0 net1
rlabel metal1 2116 6086 2116 6086 0 net10
rlabel metal1 2254 7174 2254 7174 0 net11
rlabel metal1 3496 5746 3496 5746 0 net12
rlabel metal1 6118 6766 6118 6766 0 net2
rlabel metal1 1886 3638 1886 3638 0 net3
rlabel metal1 2070 3060 2070 3060 0 net4
rlabel metal2 5198 7310 5198 7310 0 net5
rlabel metal1 5474 4114 5474 4114 0 net6
rlabel metal1 1886 4046 1886 4046 0 net7
rlabel metal1 4600 6426 4600 6426 0 net8
rlabel metal1 3818 2414 3818 2414 0 net9
rlabel metal1 6256 2550 6256 2550 0 q[0]
rlabel metal2 46 1520 46 1520 0 q[1]
rlabel metal1 6026 8058 6026 8058 0 q[2]
rlabel metal2 6486 1520 6486 1520 0 q[3]
rlabel metal3 820 3468 820 3468 0 qb[0]
rlabel metal2 5198 8194 5198 8194 0 qb[1]
rlabel metal2 3266 1520 3266 1520 0 qb[2]
rlabel metal1 1334 7514 1334 7514 0 qb[3]
rlabel metal1 3772 7854 3772 7854 0 rst
rlabel metal1 6946 6766 6946 6766 0 t
<< properties >>
string FIXED_BBOX 0 0 8258 10402
<< end >>
