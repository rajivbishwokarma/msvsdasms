MACRO FN_SIM
  ORIGIN 0 0 ;
  FOREIGN FN_SIM 0 0 ;
  SIZE 43.86 BY 49.56 ;
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 28.84 13.5 29.12 ;
      LAYER M2 ;
        RECT 1.12 38.08 13.5 38.36 ;
      LAYER M2 ;
        RECT 1.56 28.84 1.88 29.12 ;
      LAYER M3 ;
        RECT 1.58 28.98 1.86 38.22 ;
      LAYER M2 ;
        RECT 1.56 38.08 1.88 38.36 ;
    END
  END E
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 33.04 13.5 33.32 ;
      LAYER M2 ;
        RECT 1.12 33.88 13.5 34.16 ;
      LAYER M2 ;
        RECT 1.13 33.04 1.45 33.32 ;
      LAYER M3 ;
        RECT 1.15 33.18 1.43 34.02 ;
      LAYER M2 ;
        RECT 1.13 33.88 1.45 34.16 ;
      LAYER M2 ;
        RECT 1.12 42.28 13.5 42.56 ;
      LAYER M2 ;
        RECT 15.74 42.28 28.12 42.56 ;
      LAYER M2 ;
        RECT 15.74 41.44 28.12 41.72 ;
      LAYER M2 ;
        RECT 1.99 33.88 2.31 34.16 ;
      LAYER M3 ;
        RECT 2.01 34.02 2.29 42.42 ;
      LAYER M2 ;
        RECT 1.99 42.28 2.31 42.56 ;
      LAYER M2 ;
        RECT 13.33 42.28 15.91 42.56 ;
      LAYER M2 ;
        RECT 15.75 42.28 16.07 42.56 ;
      LAYER M3 ;
        RECT 15.77 41.58 16.05 42.42 ;
      LAYER M2 ;
        RECT 15.75 41.44 16.07 41.72 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 2.8 41.02 3.08 ;
      LAYER M2 ;
        RECT 15.74 46.48 28.12 46.76 ;
      LAYER M2 ;
        RECT 16.61 2.8 16.93 3.08 ;
      LAYER M3 ;
        RECT 16.63 2.94 16.91 46.62 ;
      LAYER M2 ;
        RECT 16.61 46.48 16.93 46.76 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 2.38 41.88 2.66 ;
      LAYER M2 ;
        RECT 30.36 46.48 42.74 46.76 ;
      LAYER M2 ;
        RECT 30.37 2.38 30.69 2.66 ;
      LAYER M3 ;
        RECT 30.39 2.52 30.67 46.62 ;
      LAYER M2 ;
        RECT 30.37 46.48 30.69 46.76 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 29.96 0.68 30.24 6.46 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 17.92 8.24 18.2 26.2 ;
      LAYER M3 ;
        RECT 35.98 35.12 36.26 41.32 ;
      LAYER M3 ;
        RECT 35.98 42.68 36.26 48.88 ;
      LAYER M3 ;
        RECT 17.92 26.04 18.2 34.86 ;
      LAYER M2 ;
        RECT 18.06 34.72 36.12 35 ;
      LAYER M3 ;
        RECT 35.98 34.86 36.26 35.28 ;
      LAYER M3 ;
        RECT 35.98 41.16 36.26 42.84 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 30.36 29.68 42.74 29.96 ;
      LAYER M2 ;
        RECT 30.36 37.24 42.74 37.52 ;
      LAYER M2 ;
        RECT 30.8 29.68 31.12 29.96 ;
      LAYER M3 ;
        RECT 30.82 29.82 31.1 37.38 ;
      LAYER M2 ;
        RECT 30.8 37.24 31.12 37.52 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 17.49 10.34 17.77 22.42 ;
      LAYER M2 ;
        RECT 1.12 46.48 13.5 46.76 ;
      LAYER M3 ;
        RECT 17.49 22.26 17.77 46.2 ;
      LAYER M2 ;
        RECT 13.76 46.06 17.63 46.34 ;
      LAYER M1 ;
        RECT 13.635 46.2 13.885 46.62 ;
      LAYER M2 ;
        RECT 13.33 46.48 13.76 46.76 ;
    END
  END F
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.74 29.68 28.12 29.96 ;
      LAYER M2 ;
        RECT 15.74 37.24 28.12 37.52 ;
      LAYER M2 ;
        RECT 15.75 29.68 16.07 29.96 ;
      LAYER M3 ;
        RECT 15.77 29.82 16.05 37.38 ;
      LAYER M2 ;
        RECT 15.75 37.24 16.07 37.52 ;
    END
  END C
  OBS 
  LAYER M3 ;
        RECT 7.6 26.72 7.88 32.92 ;
  LAYER M3 ;
        RECT 17.06 14.54 17.34 26.62 ;
  LAYER M3 ;
        RECT 7.6 26.46 7.88 26.88 ;
  LAYER M4 ;
        RECT 7.74 26.06 17.2 26.86 ;
  LAYER M3 ;
        RECT 17.06 26.275 17.34 26.645 ;
  LAYER M3 ;
        RECT 7.6 26.275 7.88 26.645 ;
  LAYER M4 ;
        RECT 7.575 26.06 7.905 26.86 ;
  LAYER M3 ;
        RECT 17.06 26.275 17.34 26.645 ;
  LAYER M4 ;
        RECT 17.035 26.06 17.365 26.86 ;
  LAYER M3 ;
        RECT 7.6 26.275 7.88 26.645 ;
  LAYER M4 ;
        RECT 7.575 26.06 7.905 26.86 ;
  LAYER M3 ;
        RECT 17.06 26.275 17.34 26.645 ;
  LAYER M4 ;
        RECT 17.035 26.06 17.365 26.86 ;
  LAYER M3 ;
        RECT 7.6 34.28 7.88 40.48 ;
  LAYER M3 ;
        RECT 7.6 42.68 7.88 48.88 ;
  LAYER M2 ;
        RECT 15.74 33.88 28.12 34.16 ;
  LAYER M2 ;
        RECT 30.36 33.88 42.74 34.16 ;
  LAYER M3 ;
        RECT 7.6 40.32 7.88 42.84 ;
  LAYER M3 ;
        RECT 7.6 34.02 7.88 34.44 ;
  LAYER M4 ;
        RECT 7.74 33.62 14.19 34.42 ;
  LAYER M3 ;
        RECT 14.05 33.899 14.33 34.141 ;
  LAYER M2 ;
        RECT 14.19 33.88 15.91 34.16 ;
  LAYER M2 ;
        RECT 27.95 33.88 30.53 34.16 ;
  LAYER M2 ;
        RECT 14.03 33.88 14.35 34.16 ;
  LAYER M3 ;
        RECT 14.05 33.86 14.33 34.18 ;
  LAYER M3 ;
        RECT 7.6 33.835 7.88 34.205 ;
  LAYER M4 ;
        RECT 7.575 33.62 7.905 34.42 ;
  LAYER M3 ;
        RECT 14.05 33.835 14.33 34.205 ;
  LAYER M4 ;
        RECT 14.025 33.62 14.355 34.42 ;
  LAYER M3 ;
        RECT 7.6 33.835 7.88 34.205 ;
  LAYER M4 ;
        RECT 7.575 33.62 7.905 34.42 ;
  LAYER M3 ;
        RECT 7.6 33.835 7.88 34.205 ;
  LAYER M4 ;
        RECT 7.575 33.62 7.905 34.42 ;
  LAYER M3 ;
        RECT 7.6 33.835 7.88 34.205 ;
  LAYER M4 ;
        RECT 7.575 33.62 7.905 34.42 ;
  LAYER M2 ;
        RECT 16.6 7 41.02 7.28 ;
  LAYER M3 ;
        RECT 22.22 27.56 22.5 33.76 ;
  LAYER M2 ;
        RECT 22.2 7 22.52 7.28 ;
  LAYER M3 ;
        RECT 22.22 7.14 22.5 27.72 ;
  LAYER M2 ;
        RECT 22.2 7 22.52 7.28 ;
  LAYER M3 ;
        RECT 22.22 6.98 22.5 7.3 ;
  LAYER M2 ;
        RECT 22.2 7 22.52 7.28 ;
  LAYER M3 ;
        RECT 22.22 6.98 22.5 7.3 ;
  LAYER M2 ;
        RECT 17.46 6.58 41.88 6.86 ;
  LAYER M3 ;
        RECT 35.98 27.56 36.26 33.76 ;
  LAYER M2 ;
        RECT 35.96 6.58 36.28 6.86 ;
  LAYER M3 ;
        RECT 35.98 6.72 36.26 27.72 ;
  LAYER M2 ;
        RECT 35.96 6.58 36.28 6.86 ;
  LAYER M3 ;
        RECT 35.98 6.56 36.26 6.88 ;
  LAYER M2 ;
        RECT 35.96 6.58 36.28 6.86 ;
  LAYER M3 ;
        RECT 35.98 6.56 36.26 6.88 ;
  LAYER M3 ;
        RECT 22.22 35.12 22.5 41.32 ;
  LAYER M3 ;
        RECT 22.22 42.68 22.5 48.88 ;
  LAYER M2 ;
        RECT 30.36 41.44 42.74 41.72 ;
  LAYER M2 ;
        RECT 30.36 42.28 42.74 42.56 ;
  LAYER M3 ;
        RECT 22.22 41.16 22.5 42.84 ;
  LAYER M3 ;
        RECT 22.22 41.395 22.5 41.765 ;
  LAYER M4 ;
        RECT 22.36 41.18 28.81 41.98 ;
  LAYER M3 ;
        RECT 28.67 41.459 28.95 41.701 ;
  LAYER M2 ;
        RECT 28.81 41.44 30.53 41.72 ;
  LAYER M2 ;
        RECT 30.8 41.44 31.12 41.72 ;
  LAYER M3 ;
        RECT 30.82 41.58 31.1 42.42 ;
  LAYER M2 ;
        RECT 30.8 42.28 31.12 42.56 ;
  LAYER M2 ;
        RECT 28.65 41.44 28.97 41.72 ;
  LAYER M3 ;
        RECT 28.67 41.42 28.95 41.74 ;
  LAYER M3 ;
        RECT 22.22 41.395 22.5 41.765 ;
  LAYER M4 ;
        RECT 22.195 41.18 22.525 41.98 ;
  LAYER M3 ;
        RECT 28.67 41.395 28.95 41.765 ;
  LAYER M4 ;
        RECT 28.645 41.18 28.975 41.98 ;
  LAYER M3 ;
        RECT 22.22 41.395 22.5 41.765 ;
  LAYER M4 ;
        RECT 22.195 41.18 22.525 41.98 ;
  LAYER M2 ;
        RECT 30.8 41.44 31.12 41.72 ;
  LAYER M3 ;
        RECT 30.82 41.42 31.1 41.74 ;
  LAYER M2 ;
        RECT 30.8 42.28 31.12 42.56 ;
  LAYER M3 ;
        RECT 30.82 42.26 31.1 42.58 ;
  LAYER M3 ;
        RECT 22.22 41.395 22.5 41.765 ;
  LAYER M4 ;
        RECT 22.195 41.18 22.525 41.98 ;
  LAYER M2 ;
        RECT 30.8 41.44 31.12 41.72 ;
  LAYER M3 ;
        RECT 30.82 41.42 31.1 41.74 ;
  LAYER M2 ;
        RECT 30.8 42.28 31.12 42.56 ;
  LAYER M3 ;
        RECT 30.82 42.26 31.1 42.58 ;
  LAYER M3 ;
        RECT 22.22 41.395 22.5 41.765 ;
  LAYER M4 ;
        RECT 22.195 41.18 22.525 41.98 ;
  LAYER M1 ;
        RECT 1.165 29.735 1.415 33.265 ;
  LAYER M1 ;
        RECT 1.165 28.475 1.415 29.485 ;
  LAYER M1 ;
        RECT 1.165 26.375 1.415 27.385 ;
  LAYER M1 ;
        RECT 0.735 29.735 0.985 33.265 ;
  LAYER M1 ;
        RECT 1.595 29.735 1.845 33.265 ;
  LAYER M1 ;
        RECT 2.025 29.735 2.275 33.265 ;
  LAYER M1 ;
        RECT 2.025 28.475 2.275 29.485 ;
  LAYER M1 ;
        RECT 2.025 26.375 2.275 27.385 ;
  LAYER M1 ;
        RECT 2.455 29.735 2.705 33.265 ;
  LAYER M1 ;
        RECT 2.885 29.735 3.135 33.265 ;
  LAYER M1 ;
        RECT 2.885 28.475 3.135 29.485 ;
  LAYER M1 ;
        RECT 2.885 26.375 3.135 27.385 ;
  LAYER M1 ;
        RECT 3.315 29.735 3.565 33.265 ;
  LAYER M1 ;
        RECT 3.745 29.735 3.995 33.265 ;
  LAYER M1 ;
        RECT 3.745 28.475 3.995 29.485 ;
  LAYER M1 ;
        RECT 3.745 26.375 3.995 27.385 ;
  LAYER M1 ;
        RECT 4.175 29.735 4.425 33.265 ;
  LAYER M1 ;
        RECT 4.605 29.735 4.855 33.265 ;
  LAYER M1 ;
        RECT 4.605 28.475 4.855 29.485 ;
  LAYER M1 ;
        RECT 4.605 26.375 4.855 27.385 ;
  LAYER M1 ;
        RECT 5.035 29.735 5.285 33.265 ;
  LAYER M1 ;
        RECT 5.465 29.735 5.715 33.265 ;
  LAYER M1 ;
        RECT 5.465 28.475 5.715 29.485 ;
  LAYER M1 ;
        RECT 5.465 26.375 5.715 27.385 ;
  LAYER M1 ;
        RECT 5.895 29.735 6.145 33.265 ;
  LAYER M1 ;
        RECT 6.325 29.735 6.575 33.265 ;
  LAYER M1 ;
        RECT 6.325 28.475 6.575 29.485 ;
  LAYER M1 ;
        RECT 6.325 26.375 6.575 27.385 ;
  LAYER M1 ;
        RECT 6.755 29.735 7.005 33.265 ;
  LAYER M1 ;
        RECT 7.185 29.735 7.435 33.265 ;
  LAYER M1 ;
        RECT 7.185 28.475 7.435 29.485 ;
  LAYER M1 ;
        RECT 7.185 26.375 7.435 27.385 ;
  LAYER M1 ;
        RECT 7.615 29.735 7.865 33.265 ;
  LAYER M1 ;
        RECT 8.045 29.735 8.295 33.265 ;
  LAYER M1 ;
        RECT 8.045 28.475 8.295 29.485 ;
  LAYER M1 ;
        RECT 8.045 26.375 8.295 27.385 ;
  LAYER M1 ;
        RECT 8.475 29.735 8.725 33.265 ;
  LAYER M1 ;
        RECT 8.905 29.735 9.155 33.265 ;
  LAYER M1 ;
        RECT 8.905 28.475 9.155 29.485 ;
  LAYER M1 ;
        RECT 8.905 26.375 9.155 27.385 ;
  LAYER M1 ;
        RECT 9.335 29.735 9.585 33.265 ;
  LAYER M1 ;
        RECT 9.765 29.735 10.015 33.265 ;
  LAYER M1 ;
        RECT 9.765 28.475 10.015 29.485 ;
  LAYER M1 ;
        RECT 9.765 26.375 10.015 27.385 ;
  LAYER M1 ;
        RECT 10.195 29.735 10.445 33.265 ;
  LAYER M1 ;
        RECT 10.625 29.735 10.875 33.265 ;
  LAYER M1 ;
        RECT 10.625 28.475 10.875 29.485 ;
  LAYER M1 ;
        RECT 10.625 26.375 10.875 27.385 ;
  LAYER M1 ;
        RECT 11.055 29.735 11.305 33.265 ;
  LAYER M1 ;
        RECT 11.485 29.735 11.735 33.265 ;
  LAYER M1 ;
        RECT 11.485 28.475 11.735 29.485 ;
  LAYER M1 ;
        RECT 11.485 26.375 11.735 27.385 ;
  LAYER M1 ;
        RECT 11.915 29.735 12.165 33.265 ;
  LAYER M1 ;
        RECT 12.345 29.735 12.595 33.265 ;
  LAYER M1 ;
        RECT 12.345 28.475 12.595 29.485 ;
  LAYER M1 ;
        RECT 12.345 26.375 12.595 27.385 ;
  LAYER M1 ;
        RECT 12.775 29.735 13.025 33.265 ;
  LAYER M1 ;
        RECT 13.205 29.735 13.455 33.265 ;
  LAYER M1 ;
        RECT 13.205 28.475 13.455 29.485 ;
  LAYER M1 ;
        RECT 13.205 26.375 13.455 27.385 ;
  LAYER M1 ;
        RECT 13.635 29.735 13.885 33.265 ;
  LAYER M2 ;
        RECT 0.69 32.62 13.93 32.9 ;
  LAYER M2 ;
        RECT 1.12 26.74 13.5 27.02 ;
  LAYER M2 ;
        RECT 1.12 33.04 13.5 33.32 ;
  LAYER M2 ;
        RECT 1.12 28.84 13.5 29.12 ;
  LAYER M3 ;
        RECT 7.6 26.72 7.88 32.92 ;
  LAYER M1 ;
        RECT 1.165 33.935 1.415 37.465 ;
  LAYER M1 ;
        RECT 1.165 37.715 1.415 38.725 ;
  LAYER M1 ;
        RECT 1.165 39.815 1.415 40.825 ;
  LAYER M1 ;
        RECT 0.735 33.935 0.985 37.465 ;
  LAYER M1 ;
        RECT 1.595 33.935 1.845 37.465 ;
  LAYER M1 ;
        RECT 2.025 33.935 2.275 37.465 ;
  LAYER M1 ;
        RECT 2.025 37.715 2.275 38.725 ;
  LAYER M1 ;
        RECT 2.025 39.815 2.275 40.825 ;
  LAYER M1 ;
        RECT 2.455 33.935 2.705 37.465 ;
  LAYER M1 ;
        RECT 2.885 33.935 3.135 37.465 ;
  LAYER M1 ;
        RECT 2.885 37.715 3.135 38.725 ;
  LAYER M1 ;
        RECT 2.885 39.815 3.135 40.825 ;
  LAYER M1 ;
        RECT 3.315 33.935 3.565 37.465 ;
  LAYER M1 ;
        RECT 3.745 33.935 3.995 37.465 ;
  LAYER M1 ;
        RECT 3.745 37.715 3.995 38.725 ;
  LAYER M1 ;
        RECT 3.745 39.815 3.995 40.825 ;
  LAYER M1 ;
        RECT 4.175 33.935 4.425 37.465 ;
  LAYER M1 ;
        RECT 4.605 33.935 4.855 37.465 ;
  LAYER M1 ;
        RECT 4.605 37.715 4.855 38.725 ;
  LAYER M1 ;
        RECT 4.605 39.815 4.855 40.825 ;
  LAYER M1 ;
        RECT 5.035 33.935 5.285 37.465 ;
  LAYER M1 ;
        RECT 5.465 33.935 5.715 37.465 ;
  LAYER M1 ;
        RECT 5.465 37.715 5.715 38.725 ;
  LAYER M1 ;
        RECT 5.465 39.815 5.715 40.825 ;
  LAYER M1 ;
        RECT 5.895 33.935 6.145 37.465 ;
  LAYER M1 ;
        RECT 6.325 33.935 6.575 37.465 ;
  LAYER M1 ;
        RECT 6.325 37.715 6.575 38.725 ;
  LAYER M1 ;
        RECT 6.325 39.815 6.575 40.825 ;
  LAYER M1 ;
        RECT 6.755 33.935 7.005 37.465 ;
  LAYER M1 ;
        RECT 7.185 33.935 7.435 37.465 ;
  LAYER M1 ;
        RECT 7.185 37.715 7.435 38.725 ;
  LAYER M1 ;
        RECT 7.185 39.815 7.435 40.825 ;
  LAYER M1 ;
        RECT 7.615 33.935 7.865 37.465 ;
  LAYER M1 ;
        RECT 8.045 33.935 8.295 37.465 ;
  LAYER M1 ;
        RECT 8.045 37.715 8.295 38.725 ;
  LAYER M1 ;
        RECT 8.045 39.815 8.295 40.825 ;
  LAYER M1 ;
        RECT 8.475 33.935 8.725 37.465 ;
  LAYER M1 ;
        RECT 8.905 33.935 9.155 37.465 ;
  LAYER M1 ;
        RECT 8.905 37.715 9.155 38.725 ;
  LAYER M1 ;
        RECT 8.905 39.815 9.155 40.825 ;
  LAYER M1 ;
        RECT 9.335 33.935 9.585 37.465 ;
  LAYER M1 ;
        RECT 9.765 33.935 10.015 37.465 ;
  LAYER M1 ;
        RECT 9.765 37.715 10.015 38.725 ;
  LAYER M1 ;
        RECT 9.765 39.815 10.015 40.825 ;
  LAYER M1 ;
        RECT 10.195 33.935 10.445 37.465 ;
  LAYER M1 ;
        RECT 10.625 33.935 10.875 37.465 ;
  LAYER M1 ;
        RECT 10.625 37.715 10.875 38.725 ;
  LAYER M1 ;
        RECT 10.625 39.815 10.875 40.825 ;
  LAYER M1 ;
        RECT 11.055 33.935 11.305 37.465 ;
  LAYER M1 ;
        RECT 11.485 33.935 11.735 37.465 ;
  LAYER M1 ;
        RECT 11.485 37.715 11.735 38.725 ;
  LAYER M1 ;
        RECT 11.485 39.815 11.735 40.825 ;
  LAYER M1 ;
        RECT 11.915 33.935 12.165 37.465 ;
  LAYER M1 ;
        RECT 12.345 33.935 12.595 37.465 ;
  LAYER M1 ;
        RECT 12.345 37.715 12.595 38.725 ;
  LAYER M1 ;
        RECT 12.345 39.815 12.595 40.825 ;
  LAYER M1 ;
        RECT 12.775 33.935 13.025 37.465 ;
  LAYER M1 ;
        RECT 13.205 33.935 13.455 37.465 ;
  LAYER M1 ;
        RECT 13.205 37.715 13.455 38.725 ;
  LAYER M1 ;
        RECT 13.205 39.815 13.455 40.825 ;
  LAYER M1 ;
        RECT 13.635 33.935 13.885 37.465 ;
  LAYER M2 ;
        RECT 0.69 34.3 13.93 34.58 ;
  LAYER M2 ;
        RECT 1.12 40.18 13.5 40.46 ;
  LAYER M2 ;
        RECT 1.12 33.88 13.5 34.16 ;
  LAYER M2 ;
        RECT 1.12 38.08 13.5 38.36 ;
  LAYER M3 ;
        RECT 7.6 34.28 7.88 40.48 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 18.365 3.695 18.615 7.225 ;
  LAYER M1 ;
        RECT 18.365 2.435 18.615 3.445 ;
  LAYER M1 ;
        RECT 18.365 0.335 18.615 1.345 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 20.945 3.695 21.195 7.225 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 20.945 0.335 21.195 1.345 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 23.525 3.695 23.775 7.225 ;
  LAYER M1 ;
        RECT 23.525 2.435 23.775 3.445 ;
  LAYER M1 ;
        RECT 23.525 0.335 23.775 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 1.345 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 1.345 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 31.265 2.435 31.515 3.445 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 1.345 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.985 2.435 33.235 3.445 ;
  LAYER M1 ;
        RECT 32.985 0.335 33.235 1.345 ;
  LAYER M1 ;
        RECT 33.415 3.695 33.665 7.225 ;
  LAYER M1 ;
        RECT 33.845 3.695 34.095 7.225 ;
  LAYER M1 ;
        RECT 33.845 2.435 34.095 3.445 ;
  LAYER M1 ;
        RECT 33.845 0.335 34.095 1.345 ;
  LAYER M1 ;
        RECT 34.275 3.695 34.525 7.225 ;
  LAYER M1 ;
        RECT 34.705 3.695 34.955 7.225 ;
  LAYER M1 ;
        RECT 34.705 2.435 34.955 3.445 ;
  LAYER M1 ;
        RECT 34.705 0.335 34.955 1.345 ;
  LAYER M1 ;
        RECT 35.135 3.695 35.385 7.225 ;
  LAYER M1 ;
        RECT 35.565 3.695 35.815 7.225 ;
  LAYER M1 ;
        RECT 35.565 2.435 35.815 3.445 ;
  LAYER M1 ;
        RECT 35.565 0.335 35.815 1.345 ;
  LAYER M1 ;
        RECT 35.995 3.695 36.245 7.225 ;
  LAYER M1 ;
        RECT 36.425 3.695 36.675 7.225 ;
  LAYER M1 ;
        RECT 36.425 2.435 36.675 3.445 ;
  LAYER M1 ;
        RECT 36.425 0.335 36.675 1.345 ;
  LAYER M1 ;
        RECT 36.855 3.695 37.105 7.225 ;
  LAYER M1 ;
        RECT 37.285 3.695 37.535 7.225 ;
  LAYER M1 ;
        RECT 37.285 2.435 37.535 3.445 ;
  LAYER M1 ;
        RECT 37.285 0.335 37.535 1.345 ;
  LAYER M1 ;
        RECT 37.715 3.695 37.965 7.225 ;
  LAYER M1 ;
        RECT 38.145 3.695 38.395 7.225 ;
  LAYER M1 ;
        RECT 38.145 2.435 38.395 3.445 ;
  LAYER M1 ;
        RECT 38.145 0.335 38.395 1.345 ;
  LAYER M1 ;
        RECT 38.575 3.695 38.825 7.225 ;
  LAYER M1 ;
        RECT 39.005 3.695 39.255 7.225 ;
  LAYER M1 ;
        RECT 39.005 2.435 39.255 3.445 ;
  LAYER M1 ;
        RECT 39.005 0.335 39.255 1.345 ;
  LAYER M1 ;
        RECT 39.435 3.695 39.685 7.225 ;
  LAYER M1 ;
        RECT 39.865 3.695 40.115 7.225 ;
  LAYER M1 ;
        RECT 39.865 2.435 40.115 3.445 ;
  LAYER M1 ;
        RECT 39.865 0.335 40.115 1.345 ;
  LAYER M1 ;
        RECT 40.295 3.695 40.545 7.225 ;
  LAYER M1 ;
        RECT 40.725 3.695 40.975 7.225 ;
  LAYER M1 ;
        RECT 40.725 2.435 40.975 3.445 ;
  LAYER M1 ;
        RECT 40.725 0.335 40.975 1.345 ;
  LAYER M1 ;
        RECT 41.155 3.695 41.405 7.225 ;
  LAYER M1 ;
        RECT 41.585 3.695 41.835 7.225 ;
  LAYER M1 ;
        RECT 41.585 2.435 41.835 3.445 ;
  LAYER M1 ;
        RECT 41.585 0.335 41.835 1.345 ;
  LAYER M1 ;
        RECT 42.015 3.695 42.265 7.225 ;
  LAYER M2 ;
        RECT 16.17 6.16 42.31 6.44 ;
  LAYER M2 ;
        RECT 16.6 0.7 41.88 0.98 ;
  LAYER M2 ;
        RECT 16.6 7 41.02 7.28 ;
  LAYER M2 ;
        RECT 17.46 6.58 41.88 6.86 ;
  LAYER M2 ;
        RECT 16.6 2.8 41.02 3.08 ;
  LAYER M2 ;
        RECT 17.46 2.38 41.88 2.66 ;
  LAYER M3 ;
        RECT 29.96 0.68 30.24 6.46 ;
  LAYER M1 ;
        RECT 42.445 42.335 42.695 45.865 ;
  LAYER M1 ;
        RECT 42.445 46.115 42.695 47.125 ;
  LAYER M1 ;
        RECT 42.445 48.215 42.695 49.225 ;
  LAYER M1 ;
        RECT 42.875 42.335 43.125 45.865 ;
  LAYER M1 ;
        RECT 42.015 42.335 42.265 45.865 ;
  LAYER M1 ;
        RECT 41.585 42.335 41.835 45.865 ;
  LAYER M1 ;
        RECT 41.585 46.115 41.835 47.125 ;
  LAYER M1 ;
        RECT 41.585 48.215 41.835 49.225 ;
  LAYER M1 ;
        RECT 41.155 42.335 41.405 45.865 ;
  LAYER M1 ;
        RECT 40.725 42.335 40.975 45.865 ;
  LAYER M1 ;
        RECT 40.725 46.115 40.975 47.125 ;
  LAYER M1 ;
        RECT 40.725 48.215 40.975 49.225 ;
  LAYER M1 ;
        RECT 40.295 42.335 40.545 45.865 ;
  LAYER M1 ;
        RECT 39.865 42.335 40.115 45.865 ;
  LAYER M1 ;
        RECT 39.865 46.115 40.115 47.125 ;
  LAYER M1 ;
        RECT 39.865 48.215 40.115 49.225 ;
  LAYER M1 ;
        RECT 39.435 42.335 39.685 45.865 ;
  LAYER M1 ;
        RECT 39.005 42.335 39.255 45.865 ;
  LAYER M1 ;
        RECT 39.005 46.115 39.255 47.125 ;
  LAYER M1 ;
        RECT 39.005 48.215 39.255 49.225 ;
  LAYER M1 ;
        RECT 38.575 42.335 38.825 45.865 ;
  LAYER M1 ;
        RECT 38.145 42.335 38.395 45.865 ;
  LAYER M1 ;
        RECT 38.145 46.115 38.395 47.125 ;
  LAYER M1 ;
        RECT 38.145 48.215 38.395 49.225 ;
  LAYER M1 ;
        RECT 37.715 42.335 37.965 45.865 ;
  LAYER M1 ;
        RECT 37.285 42.335 37.535 45.865 ;
  LAYER M1 ;
        RECT 37.285 46.115 37.535 47.125 ;
  LAYER M1 ;
        RECT 37.285 48.215 37.535 49.225 ;
  LAYER M1 ;
        RECT 36.855 42.335 37.105 45.865 ;
  LAYER M1 ;
        RECT 36.425 42.335 36.675 45.865 ;
  LAYER M1 ;
        RECT 36.425 46.115 36.675 47.125 ;
  LAYER M1 ;
        RECT 36.425 48.215 36.675 49.225 ;
  LAYER M1 ;
        RECT 35.995 42.335 36.245 45.865 ;
  LAYER M1 ;
        RECT 35.565 42.335 35.815 45.865 ;
  LAYER M1 ;
        RECT 35.565 46.115 35.815 47.125 ;
  LAYER M1 ;
        RECT 35.565 48.215 35.815 49.225 ;
  LAYER M1 ;
        RECT 35.135 42.335 35.385 45.865 ;
  LAYER M1 ;
        RECT 34.705 42.335 34.955 45.865 ;
  LAYER M1 ;
        RECT 34.705 46.115 34.955 47.125 ;
  LAYER M1 ;
        RECT 34.705 48.215 34.955 49.225 ;
  LAYER M1 ;
        RECT 34.275 42.335 34.525 45.865 ;
  LAYER M1 ;
        RECT 33.845 42.335 34.095 45.865 ;
  LAYER M1 ;
        RECT 33.845 46.115 34.095 47.125 ;
  LAYER M1 ;
        RECT 33.845 48.215 34.095 49.225 ;
  LAYER M1 ;
        RECT 33.415 42.335 33.665 45.865 ;
  LAYER M1 ;
        RECT 32.985 42.335 33.235 45.865 ;
  LAYER M1 ;
        RECT 32.985 46.115 33.235 47.125 ;
  LAYER M1 ;
        RECT 32.985 48.215 33.235 49.225 ;
  LAYER M1 ;
        RECT 32.555 42.335 32.805 45.865 ;
  LAYER M1 ;
        RECT 32.125 42.335 32.375 45.865 ;
  LAYER M1 ;
        RECT 32.125 46.115 32.375 47.125 ;
  LAYER M1 ;
        RECT 32.125 48.215 32.375 49.225 ;
  LAYER M1 ;
        RECT 31.695 42.335 31.945 45.865 ;
  LAYER M1 ;
        RECT 31.265 42.335 31.515 45.865 ;
  LAYER M1 ;
        RECT 31.265 46.115 31.515 47.125 ;
  LAYER M1 ;
        RECT 31.265 48.215 31.515 49.225 ;
  LAYER M1 ;
        RECT 30.835 42.335 31.085 45.865 ;
  LAYER M1 ;
        RECT 30.405 42.335 30.655 45.865 ;
  LAYER M1 ;
        RECT 30.405 46.115 30.655 47.125 ;
  LAYER M1 ;
        RECT 30.405 48.215 30.655 49.225 ;
  LAYER M1 ;
        RECT 29.975 42.335 30.225 45.865 ;
  LAYER M2 ;
        RECT 29.93 42.7 43.17 42.98 ;
  LAYER M2 ;
        RECT 30.36 48.58 42.74 48.86 ;
  LAYER M2 ;
        RECT 30.36 42.28 42.74 42.56 ;
  LAYER M2 ;
        RECT 30.36 46.48 42.74 46.76 ;
  LAYER M3 ;
        RECT 35.98 42.68 36.26 48.88 ;
  LAYER M1 ;
        RECT 42.445 38.135 42.695 41.665 ;
  LAYER M1 ;
        RECT 42.445 36.875 42.695 37.885 ;
  LAYER M1 ;
        RECT 42.445 34.775 42.695 35.785 ;
  LAYER M1 ;
        RECT 42.875 38.135 43.125 41.665 ;
  LAYER M1 ;
        RECT 42.015 38.135 42.265 41.665 ;
  LAYER M1 ;
        RECT 41.585 38.135 41.835 41.665 ;
  LAYER M1 ;
        RECT 41.585 36.875 41.835 37.885 ;
  LAYER M1 ;
        RECT 41.585 34.775 41.835 35.785 ;
  LAYER M1 ;
        RECT 41.155 38.135 41.405 41.665 ;
  LAYER M1 ;
        RECT 40.725 38.135 40.975 41.665 ;
  LAYER M1 ;
        RECT 40.725 36.875 40.975 37.885 ;
  LAYER M1 ;
        RECT 40.725 34.775 40.975 35.785 ;
  LAYER M1 ;
        RECT 40.295 38.135 40.545 41.665 ;
  LAYER M1 ;
        RECT 39.865 38.135 40.115 41.665 ;
  LAYER M1 ;
        RECT 39.865 36.875 40.115 37.885 ;
  LAYER M1 ;
        RECT 39.865 34.775 40.115 35.785 ;
  LAYER M1 ;
        RECT 39.435 38.135 39.685 41.665 ;
  LAYER M1 ;
        RECT 39.005 38.135 39.255 41.665 ;
  LAYER M1 ;
        RECT 39.005 36.875 39.255 37.885 ;
  LAYER M1 ;
        RECT 39.005 34.775 39.255 35.785 ;
  LAYER M1 ;
        RECT 38.575 38.135 38.825 41.665 ;
  LAYER M1 ;
        RECT 38.145 38.135 38.395 41.665 ;
  LAYER M1 ;
        RECT 38.145 36.875 38.395 37.885 ;
  LAYER M1 ;
        RECT 38.145 34.775 38.395 35.785 ;
  LAYER M1 ;
        RECT 37.715 38.135 37.965 41.665 ;
  LAYER M1 ;
        RECT 37.285 38.135 37.535 41.665 ;
  LAYER M1 ;
        RECT 37.285 36.875 37.535 37.885 ;
  LAYER M1 ;
        RECT 37.285 34.775 37.535 35.785 ;
  LAYER M1 ;
        RECT 36.855 38.135 37.105 41.665 ;
  LAYER M1 ;
        RECT 36.425 38.135 36.675 41.665 ;
  LAYER M1 ;
        RECT 36.425 36.875 36.675 37.885 ;
  LAYER M1 ;
        RECT 36.425 34.775 36.675 35.785 ;
  LAYER M1 ;
        RECT 35.995 38.135 36.245 41.665 ;
  LAYER M1 ;
        RECT 35.565 38.135 35.815 41.665 ;
  LAYER M1 ;
        RECT 35.565 36.875 35.815 37.885 ;
  LAYER M1 ;
        RECT 35.565 34.775 35.815 35.785 ;
  LAYER M1 ;
        RECT 35.135 38.135 35.385 41.665 ;
  LAYER M1 ;
        RECT 34.705 38.135 34.955 41.665 ;
  LAYER M1 ;
        RECT 34.705 36.875 34.955 37.885 ;
  LAYER M1 ;
        RECT 34.705 34.775 34.955 35.785 ;
  LAYER M1 ;
        RECT 34.275 38.135 34.525 41.665 ;
  LAYER M1 ;
        RECT 33.845 38.135 34.095 41.665 ;
  LAYER M1 ;
        RECT 33.845 36.875 34.095 37.885 ;
  LAYER M1 ;
        RECT 33.845 34.775 34.095 35.785 ;
  LAYER M1 ;
        RECT 33.415 38.135 33.665 41.665 ;
  LAYER M1 ;
        RECT 32.985 38.135 33.235 41.665 ;
  LAYER M1 ;
        RECT 32.985 36.875 33.235 37.885 ;
  LAYER M1 ;
        RECT 32.985 34.775 33.235 35.785 ;
  LAYER M1 ;
        RECT 32.555 38.135 32.805 41.665 ;
  LAYER M1 ;
        RECT 32.125 38.135 32.375 41.665 ;
  LAYER M1 ;
        RECT 32.125 36.875 32.375 37.885 ;
  LAYER M1 ;
        RECT 32.125 34.775 32.375 35.785 ;
  LAYER M1 ;
        RECT 31.695 38.135 31.945 41.665 ;
  LAYER M1 ;
        RECT 31.265 38.135 31.515 41.665 ;
  LAYER M1 ;
        RECT 31.265 36.875 31.515 37.885 ;
  LAYER M1 ;
        RECT 31.265 34.775 31.515 35.785 ;
  LAYER M1 ;
        RECT 30.835 38.135 31.085 41.665 ;
  LAYER M1 ;
        RECT 30.405 38.135 30.655 41.665 ;
  LAYER M1 ;
        RECT 30.405 36.875 30.655 37.885 ;
  LAYER M1 ;
        RECT 30.405 34.775 30.655 35.785 ;
  LAYER M1 ;
        RECT 29.975 38.135 30.225 41.665 ;
  LAYER M2 ;
        RECT 29.93 41.02 43.17 41.3 ;
  LAYER M2 ;
        RECT 30.36 35.14 42.74 35.42 ;
  LAYER M2 ;
        RECT 30.36 41.44 42.74 41.72 ;
  LAYER M2 ;
        RECT 30.36 37.24 42.74 37.52 ;
  LAYER M3 ;
        RECT 35.98 35.12 36.26 41.32 ;
  LAYER M1 ;
        RECT 15.785 23.015 16.035 26.545 ;
  LAYER M1 ;
        RECT 15.785 21.755 16.035 22.765 ;
  LAYER M1 ;
        RECT 15.785 17.135 16.035 20.665 ;
  LAYER M1 ;
        RECT 15.785 15.875 16.035 16.885 ;
  LAYER M1 ;
        RECT 15.785 11.255 16.035 14.785 ;
  LAYER M1 ;
        RECT 15.785 9.995 16.035 11.005 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 8.905 ;
  LAYER M1 ;
        RECT 15.355 23.015 15.605 26.545 ;
  LAYER M1 ;
        RECT 15.355 17.135 15.605 20.665 ;
  LAYER M1 ;
        RECT 15.355 11.255 15.605 14.785 ;
  LAYER M1 ;
        RECT 16.215 23.015 16.465 26.545 ;
  LAYER M1 ;
        RECT 16.215 17.135 16.465 20.665 ;
  LAYER M1 ;
        RECT 16.215 11.255 16.465 14.785 ;
  LAYER M1 ;
        RECT 16.645 23.015 16.895 26.545 ;
  LAYER M1 ;
        RECT 16.645 21.755 16.895 22.765 ;
  LAYER M1 ;
        RECT 16.645 17.135 16.895 20.665 ;
  LAYER M1 ;
        RECT 16.645 15.875 16.895 16.885 ;
  LAYER M1 ;
        RECT 16.645 11.255 16.895 14.785 ;
  LAYER M1 ;
        RECT 16.645 9.995 16.895 11.005 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 8.905 ;
  LAYER M1 ;
        RECT 17.075 23.015 17.325 26.545 ;
  LAYER M1 ;
        RECT 17.075 17.135 17.325 20.665 ;
  LAYER M1 ;
        RECT 17.075 11.255 17.325 14.785 ;
  LAYER M1 ;
        RECT 17.505 23.015 17.755 26.545 ;
  LAYER M1 ;
        RECT 17.505 21.755 17.755 22.765 ;
  LAYER M1 ;
        RECT 17.505 17.135 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.505 15.875 17.755 16.885 ;
  LAYER M1 ;
        RECT 17.505 11.255 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.505 9.995 17.755 11.005 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 8.905 ;
  LAYER M1 ;
        RECT 17.935 23.015 18.185 26.545 ;
  LAYER M1 ;
        RECT 17.935 17.135 18.185 20.665 ;
  LAYER M1 ;
        RECT 17.935 11.255 18.185 14.785 ;
  LAYER M1 ;
        RECT 18.365 23.015 18.615 26.545 ;
  LAYER M1 ;
        RECT 18.365 21.755 18.615 22.765 ;
  LAYER M1 ;
        RECT 18.365 17.135 18.615 20.665 ;
  LAYER M1 ;
        RECT 18.365 15.875 18.615 16.885 ;
  LAYER M1 ;
        RECT 18.365 11.255 18.615 14.785 ;
  LAYER M1 ;
        RECT 18.365 9.995 18.615 11.005 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 8.905 ;
  LAYER M1 ;
        RECT 18.795 23.015 19.045 26.545 ;
  LAYER M1 ;
        RECT 18.795 17.135 19.045 20.665 ;
  LAYER M1 ;
        RECT 18.795 11.255 19.045 14.785 ;
  LAYER M1 ;
        RECT 19.225 23.015 19.475 26.545 ;
  LAYER M1 ;
        RECT 19.225 21.755 19.475 22.765 ;
  LAYER M1 ;
        RECT 19.225 17.135 19.475 20.665 ;
  LAYER M1 ;
        RECT 19.225 15.875 19.475 16.885 ;
  LAYER M1 ;
        RECT 19.225 11.255 19.475 14.785 ;
  LAYER M1 ;
        RECT 19.225 9.995 19.475 11.005 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 8.905 ;
  LAYER M1 ;
        RECT 19.655 23.015 19.905 26.545 ;
  LAYER M1 ;
        RECT 19.655 17.135 19.905 20.665 ;
  LAYER M1 ;
        RECT 19.655 11.255 19.905 14.785 ;
  LAYER M2 ;
        RECT 15.74 26.32 19.52 26.6 ;
  LAYER M2 ;
        RECT 15.74 22.12 19.52 22.4 ;
  LAYER M2 ;
        RECT 15.31 25.9 19.95 26.18 ;
  LAYER M2 ;
        RECT 15.74 20.44 19.52 20.72 ;
  LAYER M2 ;
        RECT 15.74 16.24 19.52 16.52 ;
  LAYER M2 ;
        RECT 15.31 20.02 19.95 20.3 ;
  LAYER M2 ;
        RECT 15.74 14.56 19.52 14.84 ;
  LAYER M2 ;
        RECT 15.74 10.36 19.52 10.64 ;
  LAYER M2 ;
        RECT 15.31 14.14 19.95 14.42 ;
  LAYER M2 ;
        RECT 15.74 8.26 19.52 8.54 ;
  LAYER M3 ;
        RECT 17.06 14.54 17.34 26.62 ;
  LAYER M3 ;
        RECT 17.49 10.34 17.77 22.42 ;
  LAYER M3 ;
        RECT 17.92 8.24 18.2 26.2 ;
  LAYER M1 ;
        RECT 15.785 42.335 16.035 45.865 ;
  LAYER M1 ;
        RECT 15.785 46.115 16.035 47.125 ;
  LAYER M1 ;
        RECT 15.785 48.215 16.035 49.225 ;
  LAYER M1 ;
        RECT 15.355 42.335 15.605 45.865 ;
  LAYER M1 ;
        RECT 16.215 42.335 16.465 45.865 ;
  LAYER M1 ;
        RECT 16.645 42.335 16.895 45.865 ;
  LAYER M1 ;
        RECT 16.645 46.115 16.895 47.125 ;
  LAYER M1 ;
        RECT 16.645 48.215 16.895 49.225 ;
  LAYER M1 ;
        RECT 17.075 42.335 17.325 45.865 ;
  LAYER M1 ;
        RECT 17.505 42.335 17.755 45.865 ;
  LAYER M1 ;
        RECT 17.505 46.115 17.755 47.125 ;
  LAYER M1 ;
        RECT 17.505 48.215 17.755 49.225 ;
  LAYER M1 ;
        RECT 17.935 42.335 18.185 45.865 ;
  LAYER M1 ;
        RECT 18.365 42.335 18.615 45.865 ;
  LAYER M1 ;
        RECT 18.365 46.115 18.615 47.125 ;
  LAYER M1 ;
        RECT 18.365 48.215 18.615 49.225 ;
  LAYER M1 ;
        RECT 18.795 42.335 19.045 45.865 ;
  LAYER M1 ;
        RECT 19.225 42.335 19.475 45.865 ;
  LAYER M1 ;
        RECT 19.225 46.115 19.475 47.125 ;
  LAYER M1 ;
        RECT 19.225 48.215 19.475 49.225 ;
  LAYER M1 ;
        RECT 19.655 42.335 19.905 45.865 ;
  LAYER M1 ;
        RECT 20.085 42.335 20.335 45.865 ;
  LAYER M1 ;
        RECT 20.085 46.115 20.335 47.125 ;
  LAYER M1 ;
        RECT 20.085 48.215 20.335 49.225 ;
  LAYER M1 ;
        RECT 20.515 42.335 20.765 45.865 ;
  LAYER M1 ;
        RECT 20.945 42.335 21.195 45.865 ;
  LAYER M1 ;
        RECT 20.945 46.115 21.195 47.125 ;
  LAYER M1 ;
        RECT 20.945 48.215 21.195 49.225 ;
  LAYER M1 ;
        RECT 21.375 42.335 21.625 45.865 ;
  LAYER M1 ;
        RECT 21.805 42.335 22.055 45.865 ;
  LAYER M1 ;
        RECT 21.805 46.115 22.055 47.125 ;
  LAYER M1 ;
        RECT 21.805 48.215 22.055 49.225 ;
  LAYER M1 ;
        RECT 22.235 42.335 22.485 45.865 ;
  LAYER M1 ;
        RECT 22.665 42.335 22.915 45.865 ;
  LAYER M1 ;
        RECT 22.665 46.115 22.915 47.125 ;
  LAYER M1 ;
        RECT 22.665 48.215 22.915 49.225 ;
  LAYER M1 ;
        RECT 23.095 42.335 23.345 45.865 ;
  LAYER M1 ;
        RECT 23.525 42.335 23.775 45.865 ;
  LAYER M1 ;
        RECT 23.525 46.115 23.775 47.125 ;
  LAYER M1 ;
        RECT 23.525 48.215 23.775 49.225 ;
  LAYER M1 ;
        RECT 23.955 42.335 24.205 45.865 ;
  LAYER M1 ;
        RECT 24.385 42.335 24.635 45.865 ;
  LAYER M1 ;
        RECT 24.385 46.115 24.635 47.125 ;
  LAYER M1 ;
        RECT 24.385 48.215 24.635 49.225 ;
  LAYER M1 ;
        RECT 24.815 42.335 25.065 45.865 ;
  LAYER M1 ;
        RECT 25.245 42.335 25.495 45.865 ;
  LAYER M1 ;
        RECT 25.245 46.115 25.495 47.125 ;
  LAYER M1 ;
        RECT 25.245 48.215 25.495 49.225 ;
  LAYER M1 ;
        RECT 25.675 42.335 25.925 45.865 ;
  LAYER M1 ;
        RECT 26.105 42.335 26.355 45.865 ;
  LAYER M1 ;
        RECT 26.105 46.115 26.355 47.125 ;
  LAYER M1 ;
        RECT 26.105 48.215 26.355 49.225 ;
  LAYER M1 ;
        RECT 26.535 42.335 26.785 45.865 ;
  LAYER M1 ;
        RECT 26.965 42.335 27.215 45.865 ;
  LAYER M1 ;
        RECT 26.965 46.115 27.215 47.125 ;
  LAYER M1 ;
        RECT 26.965 48.215 27.215 49.225 ;
  LAYER M1 ;
        RECT 27.395 42.335 27.645 45.865 ;
  LAYER M1 ;
        RECT 27.825 42.335 28.075 45.865 ;
  LAYER M1 ;
        RECT 27.825 46.115 28.075 47.125 ;
  LAYER M1 ;
        RECT 27.825 48.215 28.075 49.225 ;
  LAYER M1 ;
        RECT 28.255 42.335 28.505 45.865 ;
  LAYER M2 ;
        RECT 15.31 42.7 28.55 42.98 ;
  LAYER M2 ;
        RECT 15.74 48.58 28.12 48.86 ;
  LAYER M2 ;
        RECT 15.74 42.28 28.12 42.56 ;
  LAYER M2 ;
        RECT 15.74 46.48 28.12 46.76 ;
  LAYER M3 ;
        RECT 22.22 42.68 22.5 48.88 ;
  LAYER M1 ;
        RECT 15.785 38.135 16.035 41.665 ;
  LAYER M1 ;
        RECT 15.785 36.875 16.035 37.885 ;
  LAYER M1 ;
        RECT 15.785 34.775 16.035 35.785 ;
  LAYER M1 ;
        RECT 15.355 38.135 15.605 41.665 ;
  LAYER M1 ;
        RECT 16.215 38.135 16.465 41.665 ;
  LAYER M1 ;
        RECT 16.645 38.135 16.895 41.665 ;
  LAYER M1 ;
        RECT 16.645 36.875 16.895 37.885 ;
  LAYER M1 ;
        RECT 16.645 34.775 16.895 35.785 ;
  LAYER M1 ;
        RECT 17.075 38.135 17.325 41.665 ;
  LAYER M1 ;
        RECT 17.505 38.135 17.755 41.665 ;
  LAYER M1 ;
        RECT 17.505 36.875 17.755 37.885 ;
  LAYER M1 ;
        RECT 17.505 34.775 17.755 35.785 ;
  LAYER M1 ;
        RECT 17.935 38.135 18.185 41.665 ;
  LAYER M1 ;
        RECT 18.365 38.135 18.615 41.665 ;
  LAYER M1 ;
        RECT 18.365 36.875 18.615 37.885 ;
  LAYER M1 ;
        RECT 18.365 34.775 18.615 35.785 ;
  LAYER M1 ;
        RECT 18.795 38.135 19.045 41.665 ;
  LAYER M1 ;
        RECT 19.225 38.135 19.475 41.665 ;
  LAYER M1 ;
        RECT 19.225 36.875 19.475 37.885 ;
  LAYER M1 ;
        RECT 19.225 34.775 19.475 35.785 ;
  LAYER M1 ;
        RECT 19.655 38.135 19.905 41.665 ;
  LAYER M1 ;
        RECT 20.085 38.135 20.335 41.665 ;
  LAYER M1 ;
        RECT 20.085 36.875 20.335 37.885 ;
  LAYER M1 ;
        RECT 20.085 34.775 20.335 35.785 ;
  LAYER M1 ;
        RECT 20.515 38.135 20.765 41.665 ;
  LAYER M1 ;
        RECT 20.945 38.135 21.195 41.665 ;
  LAYER M1 ;
        RECT 20.945 36.875 21.195 37.885 ;
  LAYER M1 ;
        RECT 20.945 34.775 21.195 35.785 ;
  LAYER M1 ;
        RECT 21.375 38.135 21.625 41.665 ;
  LAYER M1 ;
        RECT 21.805 38.135 22.055 41.665 ;
  LAYER M1 ;
        RECT 21.805 36.875 22.055 37.885 ;
  LAYER M1 ;
        RECT 21.805 34.775 22.055 35.785 ;
  LAYER M1 ;
        RECT 22.235 38.135 22.485 41.665 ;
  LAYER M1 ;
        RECT 22.665 38.135 22.915 41.665 ;
  LAYER M1 ;
        RECT 22.665 36.875 22.915 37.885 ;
  LAYER M1 ;
        RECT 22.665 34.775 22.915 35.785 ;
  LAYER M1 ;
        RECT 23.095 38.135 23.345 41.665 ;
  LAYER M1 ;
        RECT 23.525 38.135 23.775 41.665 ;
  LAYER M1 ;
        RECT 23.525 36.875 23.775 37.885 ;
  LAYER M1 ;
        RECT 23.525 34.775 23.775 35.785 ;
  LAYER M1 ;
        RECT 23.955 38.135 24.205 41.665 ;
  LAYER M1 ;
        RECT 24.385 38.135 24.635 41.665 ;
  LAYER M1 ;
        RECT 24.385 36.875 24.635 37.885 ;
  LAYER M1 ;
        RECT 24.385 34.775 24.635 35.785 ;
  LAYER M1 ;
        RECT 24.815 38.135 25.065 41.665 ;
  LAYER M1 ;
        RECT 25.245 38.135 25.495 41.665 ;
  LAYER M1 ;
        RECT 25.245 36.875 25.495 37.885 ;
  LAYER M1 ;
        RECT 25.245 34.775 25.495 35.785 ;
  LAYER M1 ;
        RECT 25.675 38.135 25.925 41.665 ;
  LAYER M1 ;
        RECT 26.105 38.135 26.355 41.665 ;
  LAYER M1 ;
        RECT 26.105 36.875 26.355 37.885 ;
  LAYER M1 ;
        RECT 26.105 34.775 26.355 35.785 ;
  LAYER M1 ;
        RECT 26.535 38.135 26.785 41.665 ;
  LAYER M1 ;
        RECT 26.965 38.135 27.215 41.665 ;
  LAYER M1 ;
        RECT 26.965 36.875 27.215 37.885 ;
  LAYER M1 ;
        RECT 26.965 34.775 27.215 35.785 ;
  LAYER M1 ;
        RECT 27.395 38.135 27.645 41.665 ;
  LAYER M1 ;
        RECT 27.825 38.135 28.075 41.665 ;
  LAYER M1 ;
        RECT 27.825 36.875 28.075 37.885 ;
  LAYER M1 ;
        RECT 27.825 34.775 28.075 35.785 ;
  LAYER M1 ;
        RECT 28.255 38.135 28.505 41.665 ;
  LAYER M2 ;
        RECT 15.31 41.02 28.55 41.3 ;
  LAYER M2 ;
        RECT 15.74 35.14 28.12 35.42 ;
  LAYER M2 ;
        RECT 15.74 41.44 28.12 41.72 ;
  LAYER M2 ;
        RECT 15.74 37.24 28.12 37.52 ;
  LAYER M3 ;
        RECT 22.22 35.12 22.5 41.32 ;
  LAYER M1 ;
        RECT 15.785 30.575 16.035 34.105 ;
  LAYER M1 ;
        RECT 15.785 29.315 16.035 30.325 ;
  LAYER M1 ;
        RECT 15.785 27.215 16.035 28.225 ;
  LAYER M1 ;
        RECT 15.355 30.575 15.605 34.105 ;
  LAYER M1 ;
        RECT 16.215 30.575 16.465 34.105 ;
  LAYER M1 ;
        RECT 16.645 30.575 16.895 34.105 ;
  LAYER M1 ;
        RECT 16.645 29.315 16.895 30.325 ;
  LAYER M1 ;
        RECT 16.645 27.215 16.895 28.225 ;
  LAYER M1 ;
        RECT 17.075 30.575 17.325 34.105 ;
  LAYER M1 ;
        RECT 17.505 30.575 17.755 34.105 ;
  LAYER M1 ;
        RECT 17.505 29.315 17.755 30.325 ;
  LAYER M1 ;
        RECT 17.505 27.215 17.755 28.225 ;
  LAYER M1 ;
        RECT 17.935 30.575 18.185 34.105 ;
  LAYER M1 ;
        RECT 18.365 30.575 18.615 34.105 ;
  LAYER M1 ;
        RECT 18.365 29.315 18.615 30.325 ;
  LAYER M1 ;
        RECT 18.365 27.215 18.615 28.225 ;
  LAYER M1 ;
        RECT 18.795 30.575 19.045 34.105 ;
  LAYER M1 ;
        RECT 19.225 30.575 19.475 34.105 ;
  LAYER M1 ;
        RECT 19.225 29.315 19.475 30.325 ;
  LAYER M1 ;
        RECT 19.225 27.215 19.475 28.225 ;
  LAYER M1 ;
        RECT 19.655 30.575 19.905 34.105 ;
  LAYER M1 ;
        RECT 20.085 30.575 20.335 34.105 ;
  LAYER M1 ;
        RECT 20.085 29.315 20.335 30.325 ;
  LAYER M1 ;
        RECT 20.085 27.215 20.335 28.225 ;
  LAYER M1 ;
        RECT 20.515 30.575 20.765 34.105 ;
  LAYER M1 ;
        RECT 20.945 30.575 21.195 34.105 ;
  LAYER M1 ;
        RECT 20.945 29.315 21.195 30.325 ;
  LAYER M1 ;
        RECT 20.945 27.215 21.195 28.225 ;
  LAYER M1 ;
        RECT 21.375 30.575 21.625 34.105 ;
  LAYER M1 ;
        RECT 21.805 30.575 22.055 34.105 ;
  LAYER M1 ;
        RECT 21.805 29.315 22.055 30.325 ;
  LAYER M1 ;
        RECT 21.805 27.215 22.055 28.225 ;
  LAYER M1 ;
        RECT 22.235 30.575 22.485 34.105 ;
  LAYER M1 ;
        RECT 22.665 30.575 22.915 34.105 ;
  LAYER M1 ;
        RECT 22.665 29.315 22.915 30.325 ;
  LAYER M1 ;
        RECT 22.665 27.215 22.915 28.225 ;
  LAYER M1 ;
        RECT 23.095 30.575 23.345 34.105 ;
  LAYER M1 ;
        RECT 23.525 30.575 23.775 34.105 ;
  LAYER M1 ;
        RECT 23.525 29.315 23.775 30.325 ;
  LAYER M1 ;
        RECT 23.525 27.215 23.775 28.225 ;
  LAYER M1 ;
        RECT 23.955 30.575 24.205 34.105 ;
  LAYER M1 ;
        RECT 24.385 30.575 24.635 34.105 ;
  LAYER M1 ;
        RECT 24.385 29.315 24.635 30.325 ;
  LAYER M1 ;
        RECT 24.385 27.215 24.635 28.225 ;
  LAYER M1 ;
        RECT 24.815 30.575 25.065 34.105 ;
  LAYER M1 ;
        RECT 25.245 30.575 25.495 34.105 ;
  LAYER M1 ;
        RECT 25.245 29.315 25.495 30.325 ;
  LAYER M1 ;
        RECT 25.245 27.215 25.495 28.225 ;
  LAYER M1 ;
        RECT 25.675 30.575 25.925 34.105 ;
  LAYER M1 ;
        RECT 26.105 30.575 26.355 34.105 ;
  LAYER M1 ;
        RECT 26.105 29.315 26.355 30.325 ;
  LAYER M1 ;
        RECT 26.105 27.215 26.355 28.225 ;
  LAYER M1 ;
        RECT 26.535 30.575 26.785 34.105 ;
  LAYER M1 ;
        RECT 26.965 30.575 27.215 34.105 ;
  LAYER M1 ;
        RECT 26.965 29.315 27.215 30.325 ;
  LAYER M1 ;
        RECT 26.965 27.215 27.215 28.225 ;
  LAYER M1 ;
        RECT 27.395 30.575 27.645 34.105 ;
  LAYER M1 ;
        RECT 27.825 30.575 28.075 34.105 ;
  LAYER M1 ;
        RECT 27.825 29.315 28.075 30.325 ;
  LAYER M1 ;
        RECT 27.825 27.215 28.075 28.225 ;
  LAYER M1 ;
        RECT 28.255 30.575 28.505 34.105 ;
  LAYER M2 ;
        RECT 15.31 33.46 28.55 33.74 ;
  LAYER M2 ;
        RECT 15.74 27.58 28.12 27.86 ;
  LAYER M2 ;
        RECT 15.74 33.88 28.12 34.16 ;
  LAYER M2 ;
        RECT 15.74 29.68 28.12 29.96 ;
  LAYER M3 ;
        RECT 22.22 27.56 22.5 33.76 ;
  LAYER M1 ;
        RECT 42.445 30.575 42.695 34.105 ;
  LAYER M1 ;
        RECT 42.445 29.315 42.695 30.325 ;
  LAYER M1 ;
        RECT 42.445 27.215 42.695 28.225 ;
  LAYER M1 ;
        RECT 42.875 30.575 43.125 34.105 ;
  LAYER M1 ;
        RECT 42.015 30.575 42.265 34.105 ;
  LAYER M1 ;
        RECT 41.585 30.575 41.835 34.105 ;
  LAYER M1 ;
        RECT 41.585 29.315 41.835 30.325 ;
  LAYER M1 ;
        RECT 41.585 27.215 41.835 28.225 ;
  LAYER M1 ;
        RECT 41.155 30.575 41.405 34.105 ;
  LAYER M1 ;
        RECT 40.725 30.575 40.975 34.105 ;
  LAYER M1 ;
        RECT 40.725 29.315 40.975 30.325 ;
  LAYER M1 ;
        RECT 40.725 27.215 40.975 28.225 ;
  LAYER M1 ;
        RECT 40.295 30.575 40.545 34.105 ;
  LAYER M1 ;
        RECT 39.865 30.575 40.115 34.105 ;
  LAYER M1 ;
        RECT 39.865 29.315 40.115 30.325 ;
  LAYER M1 ;
        RECT 39.865 27.215 40.115 28.225 ;
  LAYER M1 ;
        RECT 39.435 30.575 39.685 34.105 ;
  LAYER M1 ;
        RECT 39.005 30.575 39.255 34.105 ;
  LAYER M1 ;
        RECT 39.005 29.315 39.255 30.325 ;
  LAYER M1 ;
        RECT 39.005 27.215 39.255 28.225 ;
  LAYER M1 ;
        RECT 38.575 30.575 38.825 34.105 ;
  LAYER M1 ;
        RECT 38.145 30.575 38.395 34.105 ;
  LAYER M1 ;
        RECT 38.145 29.315 38.395 30.325 ;
  LAYER M1 ;
        RECT 38.145 27.215 38.395 28.225 ;
  LAYER M1 ;
        RECT 37.715 30.575 37.965 34.105 ;
  LAYER M1 ;
        RECT 37.285 30.575 37.535 34.105 ;
  LAYER M1 ;
        RECT 37.285 29.315 37.535 30.325 ;
  LAYER M1 ;
        RECT 37.285 27.215 37.535 28.225 ;
  LAYER M1 ;
        RECT 36.855 30.575 37.105 34.105 ;
  LAYER M1 ;
        RECT 36.425 30.575 36.675 34.105 ;
  LAYER M1 ;
        RECT 36.425 29.315 36.675 30.325 ;
  LAYER M1 ;
        RECT 36.425 27.215 36.675 28.225 ;
  LAYER M1 ;
        RECT 35.995 30.575 36.245 34.105 ;
  LAYER M1 ;
        RECT 35.565 30.575 35.815 34.105 ;
  LAYER M1 ;
        RECT 35.565 29.315 35.815 30.325 ;
  LAYER M1 ;
        RECT 35.565 27.215 35.815 28.225 ;
  LAYER M1 ;
        RECT 35.135 30.575 35.385 34.105 ;
  LAYER M1 ;
        RECT 34.705 30.575 34.955 34.105 ;
  LAYER M1 ;
        RECT 34.705 29.315 34.955 30.325 ;
  LAYER M1 ;
        RECT 34.705 27.215 34.955 28.225 ;
  LAYER M1 ;
        RECT 34.275 30.575 34.525 34.105 ;
  LAYER M1 ;
        RECT 33.845 30.575 34.095 34.105 ;
  LAYER M1 ;
        RECT 33.845 29.315 34.095 30.325 ;
  LAYER M1 ;
        RECT 33.845 27.215 34.095 28.225 ;
  LAYER M1 ;
        RECT 33.415 30.575 33.665 34.105 ;
  LAYER M1 ;
        RECT 32.985 30.575 33.235 34.105 ;
  LAYER M1 ;
        RECT 32.985 29.315 33.235 30.325 ;
  LAYER M1 ;
        RECT 32.985 27.215 33.235 28.225 ;
  LAYER M1 ;
        RECT 32.555 30.575 32.805 34.105 ;
  LAYER M1 ;
        RECT 32.125 30.575 32.375 34.105 ;
  LAYER M1 ;
        RECT 32.125 29.315 32.375 30.325 ;
  LAYER M1 ;
        RECT 32.125 27.215 32.375 28.225 ;
  LAYER M1 ;
        RECT 31.695 30.575 31.945 34.105 ;
  LAYER M1 ;
        RECT 31.265 30.575 31.515 34.105 ;
  LAYER M1 ;
        RECT 31.265 29.315 31.515 30.325 ;
  LAYER M1 ;
        RECT 31.265 27.215 31.515 28.225 ;
  LAYER M1 ;
        RECT 30.835 30.575 31.085 34.105 ;
  LAYER M1 ;
        RECT 30.405 30.575 30.655 34.105 ;
  LAYER M1 ;
        RECT 30.405 29.315 30.655 30.325 ;
  LAYER M1 ;
        RECT 30.405 27.215 30.655 28.225 ;
  LAYER M1 ;
        RECT 29.975 30.575 30.225 34.105 ;
  LAYER M2 ;
        RECT 29.93 33.46 43.17 33.74 ;
  LAYER M2 ;
        RECT 30.36 27.58 42.74 27.86 ;
  LAYER M2 ;
        RECT 30.36 33.88 42.74 34.16 ;
  LAYER M2 ;
        RECT 30.36 29.68 42.74 29.96 ;
  LAYER M3 ;
        RECT 35.98 27.56 36.26 33.76 ;
  LAYER M1 ;
        RECT 1.165 42.335 1.415 45.865 ;
  LAYER M1 ;
        RECT 1.165 46.115 1.415 47.125 ;
  LAYER M1 ;
        RECT 1.165 48.215 1.415 49.225 ;
  LAYER M1 ;
        RECT 0.735 42.335 0.985 45.865 ;
  LAYER M1 ;
        RECT 1.595 42.335 1.845 45.865 ;
  LAYER M1 ;
        RECT 2.025 42.335 2.275 45.865 ;
  LAYER M1 ;
        RECT 2.025 46.115 2.275 47.125 ;
  LAYER M1 ;
        RECT 2.025 48.215 2.275 49.225 ;
  LAYER M1 ;
        RECT 2.455 42.335 2.705 45.865 ;
  LAYER M1 ;
        RECT 2.885 42.335 3.135 45.865 ;
  LAYER M1 ;
        RECT 2.885 46.115 3.135 47.125 ;
  LAYER M1 ;
        RECT 2.885 48.215 3.135 49.225 ;
  LAYER M1 ;
        RECT 3.315 42.335 3.565 45.865 ;
  LAYER M1 ;
        RECT 3.745 42.335 3.995 45.865 ;
  LAYER M1 ;
        RECT 3.745 46.115 3.995 47.125 ;
  LAYER M1 ;
        RECT 3.745 48.215 3.995 49.225 ;
  LAYER M1 ;
        RECT 4.175 42.335 4.425 45.865 ;
  LAYER M1 ;
        RECT 4.605 42.335 4.855 45.865 ;
  LAYER M1 ;
        RECT 4.605 46.115 4.855 47.125 ;
  LAYER M1 ;
        RECT 4.605 48.215 4.855 49.225 ;
  LAYER M1 ;
        RECT 5.035 42.335 5.285 45.865 ;
  LAYER M1 ;
        RECT 5.465 42.335 5.715 45.865 ;
  LAYER M1 ;
        RECT 5.465 46.115 5.715 47.125 ;
  LAYER M1 ;
        RECT 5.465 48.215 5.715 49.225 ;
  LAYER M1 ;
        RECT 5.895 42.335 6.145 45.865 ;
  LAYER M1 ;
        RECT 6.325 42.335 6.575 45.865 ;
  LAYER M1 ;
        RECT 6.325 46.115 6.575 47.125 ;
  LAYER M1 ;
        RECT 6.325 48.215 6.575 49.225 ;
  LAYER M1 ;
        RECT 6.755 42.335 7.005 45.865 ;
  LAYER M1 ;
        RECT 7.185 42.335 7.435 45.865 ;
  LAYER M1 ;
        RECT 7.185 46.115 7.435 47.125 ;
  LAYER M1 ;
        RECT 7.185 48.215 7.435 49.225 ;
  LAYER M1 ;
        RECT 7.615 42.335 7.865 45.865 ;
  LAYER M1 ;
        RECT 8.045 42.335 8.295 45.865 ;
  LAYER M1 ;
        RECT 8.045 46.115 8.295 47.125 ;
  LAYER M1 ;
        RECT 8.045 48.215 8.295 49.225 ;
  LAYER M1 ;
        RECT 8.475 42.335 8.725 45.865 ;
  LAYER M1 ;
        RECT 8.905 42.335 9.155 45.865 ;
  LAYER M1 ;
        RECT 8.905 46.115 9.155 47.125 ;
  LAYER M1 ;
        RECT 8.905 48.215 9.155 49.225 ;
  LAYER M1 ;
        RECT 9.335 42.335 9.585 45.865 ;
  LAYER M1 ;
        RECT 9.765 42.335 10.015 45.865 ;
  LAYER M1 ;
        RECT 9.765 46.115 10.015 47.125 ;
  LAYER M1 ;
        RECT 9.765 48.215 10.015 49.225 ;
  LAYER M1 ;
        RECT 10.195 42.335 10.445 45.865 ;
  LAYER M1 ;
        RECT 10.625 42.335 10.875 45.865 ;
  LAYER M1 ;
        RECT 10.625 46.115 10.875 47.125 ;
  LAYER M1 ;
        RECT 10.625 48.215 10.875 49.225 ;
  LAYER M1 ;
        RECT 11.055 42.335 11.305 45.865 ;
  LAYER M1 ;
        RECT 11.485 42.335 11.735 45.865 ;
  LAYER M1 ;
        RECT 11.485 46.115 11.735 47.125 ;
  LAYER M1 ;
        RECT 11.485 48.215 11.735 49.225 ;
  LAYER M1 ;
        RECT 11.915 42.335 12.165 45.865 ;
  LAYER M1 ;
        RECT 12.345 42.335 12.595 45.865 ;
  LAYER M1 ;
        RECT 12.345 46.115 12.595 47.125 ;
  LAYER M1 ;
        RECT 12.345 48.215 12.595 49.225 ;
  LAYER M1 ;
        RECT 12.775 42.335 13.025 45.865 ;
  LAYER M1 ;
        RECT 13.205 42.335 13.455 45.865 ;
  LAYER M1 ;
        RECT 13.205 46.115 13.455 47.125 ;
  LAYER M1 ;
        RECT 13.205 48.215 13.455 49.225 ;
  LAYER M1 ;
        RECT 13.635 42.335 13.885 45.865 ;
  LAYER M2 ;
        RECT 0.69 42.7 13.93 42.98 ;
  LAYER M2 ;
        RECT 1.12 48.58 13.5 48.86 ;
  LAYER M2 ;
        RECT 1.12 42.28 13.5 42.56 ;
  LAYER M2 ;
        RECT 1.12 46.48 13.5 46.76 ;
  LAYER M3 ;
        RECT 7.6 42.68 7.88 48.88 ;
  END 
END FN_SIM
