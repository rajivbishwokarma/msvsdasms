* SPICE3 file created from fnc.ext - technology: sky130A

.subckt fnc A C E F D B gnd vdd Fn
X0 vdd F a_190_270# vdd sky130_fd_pr__pfet_01v8 ad=1.95e+12p pd=1.19e+07u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 a_190_270# E vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n70_270# A vdd vdd sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X3 gnd F a_190_n70# Fn sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X4 vdd B a_450_270# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X5 a_190_n70# E Fn Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.5e+11p ps=5.9e+06u w=1e+06u l=150000u
X6 a_450_270# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n70_n70# A Fn Fn sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X8 gnd B a_n70_n70# Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n70_n70# D gnd Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 vdd C a_n70_270# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Fn C a_n70_n70# Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 gnd A 0.03fF
C1 A C 0.08fF
C2 a_190_270# A 0.00fF
C3 E vdd 0.07fF
C4 F vdd 0.07fF
C5 gnd vdd 0.24fF
C6 a_n70_n70# E 0.06fF
C7 C vdd 0.07fF
C8 a_190_270# vdd 0.09fF
C9 D vdd 0.07fF
C10 a_190_n70# F 0.00fF
C11 a_n70_n70# F 0.03fF
C12 gnd a_190_n70# 0.01fF
C13 a_450_270# vdd 0.04fF
C14 gnd a_n70_n70# 0.61fF
C15 a_n70_n70# C 0.05fF
C16 gnd a_n70_270# 0.00fF
C17 a_190_270# a_n70_270# 0.00fF
C18 gnd B 0.03fF
C19 a_n70_n70# D 0.03fF
C20 A vdd 0.09fF
C21 a_190_270# B 0.00fF
C22 B D 0.08fF
C23 a_n70_n70# A 0.02fF
C24 F E 0.08fF
C25 gnd E 0.02fF
C26 E C 0.08fF
C27 a_190_270# E 0.00fF
C28 gnd F 0.03fF
C29 a_190_n70# vdd 0.00fF
C30 a_190_270# F 0.00fF
C31 gnd C 0.02fF
C32 a_n70_n70# vdd 0.00fF
C33 a_n70_270# vdd 0.04fF
C34 gnd a_190_270# 0.00fF
C35 D F 0.08fF
C36 a_190_270# C 0.00fF
C37 gnd D 0.05fF
C38 B vdd 0.08fF
C39 a_190_270# D 0.00fF
C40 gnd a_450_270# 0.00fF
C41 a_190_n70# a_n70_n70# 0.03fF
C42 a_190_270# a_450_270# 0.00fF
C43 a_n70_n70# B 0.03fF
C44 gnd Fn 0.78fF
C45 B Fn 0.24fF
C46 D Fn 0.18fF
C47 F Fn 0.18fF
C48 E Fn 0.20fF
C49 C Fn 0.19fF
C50 A Fn 0.27fF
C51 vdd Fn 2.67fF
C52 a_190_n70# Fn 0.01fF **FLOATING
C53 a_n70_n70# Fn 0.14fF **FLOATING
C54 a_450_270# Fn 0.03fF **FLOATING
C55 a_190_270# Fn 0.08fF **FLOATING
C56 a_n70_270# Fn 0.02fF **FLOATING
.ends
