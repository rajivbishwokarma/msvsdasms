magic
tech sky130A
timestamp 1676090261
<< nwell >>
rect -165 100 360 270
<< nmos >>
rect -50 -35 -35 65
rect 15 -35 30 65
rect 80 -35 95 65
rect 145 -35 160 65
rect 210 -35 225 65
rect 275 -35 290 65
<< pmos >>
rect -50 135 -35 235
rect 15 135 30 235
rect 80 135 95 235
rect 145 135 160 235
rect 210 135 225 235
rect 275 135 290 235
<< ndiff >>
rect -95 55 -50 65
rect -95 30 -85 55
rect -65 30 -50 55
rect -95 0 -50 30
rect -95 -25 -85 0
rect -65 -25 -50 0
rect -95 -35 -50 -25
rect -35 55 15 65
rect -35 -25 -20 55
rect 0 -25 15 55
rect -35 -35 15 -25
rect 30 55 80 65
rect 30 30 45 55
rect 65 30 80 55
rect 30 -35 80 30
rect 95 -35 145 65
rect 160 0 210 65
rect 160 -25 175 0
rect 195 -25 210 0
rect 160 -35 210 -25
rect 225 55 275 65
rect 225 -25 240 55
rect 260 -25 275 55
rect 225 -35 275 -25
rect 290 55 340 65
rect 290 30 305 55
rect 325 30 340 55
rect 290 0 340 30
rect 290 -25 305 0
rect 325 -25 340 0
rect 290 -35 340 -25
<< pdiff >>
rect -95 225 -50 235
rect -95 200 -85 225
rect -65 200 -50 225
rect -95 170 -50 200
rect -95 145 -85 170
rect -65 145 -50 170
rect -95 135 -50 145
rect -35 135 15 235
rect 30 225 80 235
rect 30 200 45 225
rect 65 200 80 225
rect 30 135 80 200
rect 95 170 145 235
rect 95 145 110 170
rect 130 145 145 170
rect 95 135 145 145
rect 160 225 210 235
rect 160 200 175 225
rect 195 200 210 225
rect 160 135 210 200
rect 225 135 275 235
rect 290 225 340 235
rect 290 200 305 225
rect 325 200 340 225
rect 290 170 340 200
rect 290 145 305 170
rect 325 145 340 170
rect 290 135 340 145
<< ndiffc >>
rect -85 30 -65 55
rect -85 -25 -65 0
rect -20 -25 0 55
rect 45 30 65 55
rect 175 -25 195 0
rect 240 -25 260 55
rect 305 30 325 55
rect 305 -25 325 0
<< pdiffc >>
rect -85 200 -65 225
rect -85 145 -65 170
rect 45 200 65 225
rect 110 145 130 170
rect 175 200 195 225
rect 305 200 325 225
rect 305 145 325 170
<< psubdiff >>
rect -145 55 -95 65
rect -145 30 -125 55
rect -105 30 -95 55
rect -145 0 -95 30
rect -145 -25 -125 0
rect -105 -25 -95 0
rect -145 -35 -95 -25
<< nsubdiff >>
rect -145 225 -95 235
rect -145 200 -125 225
rect -105 200 -95 225
rect -145 170 -95 200
rect -145 145 -125 170
rect -105 145 -95 170
rect -145 135 -95 145
<< psubdiffcont >>
rect -125 30 -105 55
rect -125 -25 -105 0
<< nsubdiffcont >>
rect -125 200 -105 225
rect -125 145 -105 170
<< poly >>
rect -50 235 -35 250
rect 15 235 30 250
rect 80 235 95 250
rect 145 235 160 250
rect 210 235 225 250
rect 275 235 290 250
rect -50 65 -35 135
rect 15 65 30 135
rect 80 65 95 135
rect 145 65 160 135
rect 210 65 225 135
rect 275 65 290 135
rect -50 -50 -35 -35
rect 15 -50 30 -35
rect 80 -50 95 -35
rect 145 -50 160 -35
rect 210 -50 225 -35
rect 275 -50 290 -35
rect -75 -60 -35 -50
rect -75 -80 -65 -60
rect -45 -80 -35 -60
rect -75 -90 -35 -80
rect -10 -60 30 -50
rect -10 -80 0 -60
rect 20 -80 30 -60
rect -10 -90 30 -80
rect 55 -60 95 -50
rect 55 -80 65 -60
rect 85 -80 95 -60
rect 55 -90 95 -80
rect 120 -60 160 -50
rect 120 -80 130 -60
rect 150 -80 160 -60
rect 120 -90 160 -80
rect 185 -60 225 -50
rect 185 -80 195 -60
rect 215 -80 225 -60
rect 185 -90 225 -80
rect 250 -60 290 -50
rect 250 -80 260 -60
rect 280 -80 290 -60
rect 250 -90 290 -80
<< polycont >>
rect -65 -80 -45 -60
rect 0 -80 20 -60
rect 65 -80 85 -60
rect 130 -80 150 -60
rect 195 -80 215 -60
rect 260 -80 280 -60
<< locali >>
rect -135 225 -55 230
rect -135 145 -125 225
rect -105 145 -85 225
rect -65 145 -55 225
rect 35 225 75 230
rect 35 200 45 225
rect 65 200 75 225
rect 35 195 75 200
rect 165 225 205 230
rect 165 200 175 225
rect 195 200 205 225
rect 165 195 205 200
rect 295 225 335 230
rect 295 195 305 225
rect -135 140 -55 145
rect 100 170 140 175
rect 100 145 110 170
rect 130 145 140 170
rect 100 140 140 145
rect 295 145 305 175
rect 325 195 335 225
rect 325 145 335 175
rect 295 140 335 145
rect -165 90 360 110
rect -85 60 -65 90
rect 45 60 65 90
rect -135 55 -55 60
rect -135 30 -125 55
rect -105 30 -85 55
rect -65 30 -55 55
rect -135 0 -55 30
rect -135 -25 -125 0
rect -105 -25 -85 0
rect -65 -25 -55 0
rect -135 -30 -55 -25
rect -30 55 10 60
rect -30 -25 -20 55
rect 0 0 10 55
rect 35 55 75 60
rect 35 30 45 55
rect 65 30 75 55
rect 230 55 270 60
rect 230 45 240 55
rect 35 25 75 30
rect 100 25 240 45
rect 100 0 120 25
rect 0 -20 120 0
rect 165 0 205 5
rect 0 -25 10 -20
rect -30 -30 10 -25
rect 165 -25 175 0
rect 195 -25 205 0
rect 165 -30 205 -25
rect 230 -25 240 25
rect 260 -25 270 55
rect 295 55 335 60
rect 295 25 305 55
rect 230 -30 270 -25
rect 295 -25 305 5
rect 325 25 335 55
rect 325 -25 335 5
rect 295 -30 335 -25
rect -75 -60 -35 -50
rect -75 -80 -65 -60
rect -45 -80 -35 -60
rect -75 -90 -35 -80
rect -10 -60 30 -50
rect -10 -80 0 -60
rect 20 -80 30 -60
rect -10 -90 30 -80
rect 55 -60 95 -50
rect 55 -80 65 -60
rect 85 -80 95 -60
rect 55 -90 95 -80
rect 120 -60 160 -50
rect 120 -80 130 -60
rect 150 -80 160 -60
rect 120 -90 160 -80
rect 185 -60 225 -50
rect 185 -80 195 -60
rect 215 -80 225 -60
rect 185 -90 225 -80
rect 250 -60 290 -50
rect 250 -80 260 -60
rect 280 -80 290 -60
rect 250 -90 290 -80
<< viali >>
rect -125 200 -105 225
rect -125 170 -105 200
rect -125 145 -105 170
rect -85 200 -65 225
rect -85 170 -65 200
rect -85 145 -65 170
rect 45 200 65 225
rect 175 200 195 225
rect 305 200 325 225
rect 305 170 325 200
rect 305 145 325 170
rect 175 -25 195 0
rect 305 30 325 55
rect 305 0 325 30
rect 305 -25 325 0
<< metal1 >>
rect -165 225 360 230
rect -165 145 -125 225
rect -105 145 -85 225
rect -65 200 45 225
rect 65 200 175 225
rect 195 200 305 225
rect -65 145 305 200
rect 325 145 360 225
rect -165 140 360 145
rect -165 55 360 60
rect -165 0 305 55
rect -165 -25 175 0
rect 195 -25 305 0
rect 325 -25 360 55
rect -165 -30 360 -25
<< labels >>
rlabel locali -70 -70 -70 -70 1 A
port 1 n
rlabel locali -5 -70 -5 -70 1 C
port 2 n
rlabel locali 60 -70 60 -70 1 E
port 3 n
rlabel locali 125 -70 125 -70 1 F
port 4 n
rlabel locali 190 -70 190 -70 1 D
port 5 n
rlabel locali 255 -70 255 -70 1 B
port 6 n
rlabel locali 360 100 360 100 7 Fn
port 7 w
rlabel metal1 -165 185 -165 185 7 vdd
port 8 w
rlabel metal1 -165 10 -165 10 7 gnd
port 9 w
<< end >>
