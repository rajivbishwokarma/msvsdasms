* SPICE3 file created from fnc.ext - technology: sky130A

.subckt fnc A C E F D B gnd vdd Fn
X0 vdd F a_190_270# vdd sky130_fd_pr__pfet_01v8 ad=1.95e+12p pd=1.19e+07u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 a_190_270# E vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n70_270# A vdd vdd sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X3 gnd F a_190_n70# Fn sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X4 vdd B a_450_270# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X5 a_190_n70# E Fn Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.5e+11p ps=5.9e+06u w=1e+06u l=150000u
X6 a_450_270# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n70_n70# A Fn Fn sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X8 gnd B a_n70_n70# Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n70_n70# D gnd Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 vdd C a_n70_270# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Fn C a_n70_n70# Fn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 D B 0.08fF
C1 vdd a_190_270# 0.09fF
C2 a_n70_n70# vdd 0.00fF
C3 a_n70_270# gnd 0.00fF
C4 B gnd 0.03fF
C5 D vdd 0.07fF
C6 D a_190_270# 0.00fF
C7 D a_n70_n70# 0.03fF
C8 E vdd 0.07fF
C9 vdd a_190_n70# 0.00fF
C10 E a_190_270# 0.00fF
C11 E a_n70_n70# 0.06fF
C12 a_n70_n70# a_190_n70# 0.03fF
C13 vdd gnd 0.24fF
C14 a_190_270# gnd 0.00fF
C15 a_n70_n70# gnd 0.61fF
C16 vdd F 0.07fF
C17 vdd A 0.09fF
C18 F a_190_270# 0.00fF
C19 a_n70_n70# F 0.03fF
C20 A a_190_270# 0.00fF
C21 a_n70_n70# A 0.02fF
C22 D gnd 0.05fF
C23 vdd C 0.07fF
C24 C a_190_270# 0.00fF
C25 a_n70_n70# C 0.05fF
C26 vdd a_450_270# 0.04fF
C27 E gnd 0.02fF
C28 a_190_n70# gnd 0.01fF
C29 a_450_270# a_190_270# 0.00fF
C30 D F 0.08fF
C31 E F 0.08fF
C32 a_190_n70# F 0.00fF
C33 E C 0.08fF
C34 F gnd 0.03fF
C35 A gnd 0.03fF
C36 C gnd 0.02fF
C37 a_450_270# gnd 0.00fF
C38 C A 0.08fF
C39 vdd a_n70_270# 0.04fF
C40 a_n70_270# a_190_270# 0.00fF
C41 vdd B 0.08fF
C42 a_190_270# B 0.00fF
C43 a_n70_n70# B 0.03fF
C44 gnd Fn 0.78fF
C45 B Fn 0.24fF
C46 D Fn 0.18fF
C47 F Fn 0.18fF
C48 E Fn 0.20fF
C49 C Fn 0.19fF
C50 A Fn 0.27fF
C51 vdd Fn 2.67fF
C52 a_190_n70# Fn 0.01fF **FLOATING
C53 a_n70_n70# Fn 0.14fF **FLOATING
C54 a_450_270# Fn 0.03fF **FLOATING
C55 a_190_270# Fn 0.08fF **FLOATING
C56 a_n70_270# Fn 0.02fF **FLOATING
.ends
