* SPICE3 file created from RING_OSC_0.ext - technology: sky130A

.option scale=5000u

X0 li_405_1579# STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# SUB SUB sky130_fd_pr__nfet_01v8 ad=4704 pd=280 as=26712 ps=1644 w=84 l=30
X1 SUB STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# li_405_1579# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X2 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# li_663_2335# SUB SUB sky130_fd_pr__nfet_01v8 ad=4704 pd=280 as=0 ps=0 w=84 l=30
X3 SUB li_663_2335# STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X4 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# li_663_2335# m1_312_3080# m1_312_3080# sky130_fd_pr__pfet_01v8 ad=4704 pd=280 as=26712 ps=1644 w=84 l=30
X5 m1_312_3080# li_663_2335# STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# m1_312_3080# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X6 li_405_1579# STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# m1_312_3080# m1_312_3080# sky130_fd_pr__pfet_01v8 ad=4704 pd=280 as=0 ps=0 w=84 l=30
X7 m1_312_3080# STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# li_405_1579# m1_312_3080# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X8 li_663_2335# li_405_1579# m1_312_3080# m1_312_3080# sky130_fd_pr__pfet_01v8 ad=4704 pd=280 as=0 ps=0 w=84 l=30
X9 m1_312_3080# li_405_1579# li_663_2335# m1_312_3080# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X10 li_663_2335# li_405_1579# SUB SUB sky130_fd_pr__nfet_01v8 ad=4704 pd=280 as=0 ps=0 w=84 l=30
X11 SUB li_405_1579# li_663_2335# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
C0 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# VDD 0.01fF
C1 GND li_405_1579# 0.05fF
C2 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# Y 0.05fF
C3 li_663_2335# STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# 0.60fF
C4 li_663_2335# m1_312_3080# 2.26fF
C5 GND VDD 0.23fF
C6 VDD li_405_1579# 1.24fF
C7 GND Y 0.05fF
C8 li_663_2335# li_405_1579# 0.65fF
C9 VDD Y 0.31fF
C10 li_663_2335# VDD 0.55fF
C11 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# m1_312_3080# 3.00fF
C12 GND STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# 0.10fF
C13 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# li_405_1579# 0.50fF
C14 m1_312_3080# li_405_1579# 2.17fF
C15 VDD SUB 0.15fF
C16 li_405_1579# SUB 2.24fF **FLOATING
C17 STAGE2_INV_5734008_0_0_1677543509_0/li_577_571# SUB 1.17fF **FLOATING
C18 m1_312_3080# SUB 7.98fF **FLOATING
C19 li_663_2335# SUB 2.80fF **FLOATING
