MACRO FN_SIM
  ORIGIN 0 0 ;
  FOREIGN FN_SIM 0 0 ;
  SIZE 39.56 BY 33.18 ;
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.45 5.74 22.53 6.02 ;
      LAYER M2 ;
        RECT 14.45 14.98 22.53 15.26 ;
      LAYER M2 ;
        RECT 14.89 5.74 15.21 6.02 ;
      LAYER M3 ;
        RECT 14.91 5.88 15.19 15.12 ;
      LAYER M2 ;
        RECT 14.89 14.98 15.21 15.26 ;
    END
  END E
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 9.75 11.6 10.03 17.8 ;
      LAYER M2 ;
        RECT 14.45 9.94 22.53 10.22 ;
      LAYER M2 ;
        RECT 14.45 10.78 22.53 11.06 ;
      LAYER M2 ;
        RECT 14.46 9.94 14.78 10.22 ;
      LAYER M3 ;
        RECT 14.48 10.08 14.76 10.92 ;
      LAYER M2 ;
        RECT 14.46 10.78 14.78 11.06 ;
      LAYER M2 ;
        RECT 17.03 18.34 25.11 18.62 ;
      LAYER M2 ;
        RECT 27.35 18.34 35.43 18.62 ;
      LAYER M3 ;
        RECT 9.75 10.92 10.03 11.76 ;
      LAYER M2 ;
        RECT 9.89 10.78 14.62 11.06 ;
      LAYER M2 ;
        RECT 17.04 10.78 17.36 11.06 ;
      LAYER M3 ;
        RECT 17.06 10.92 17.34 18.48 ;
      LAYER M2 ;
        RECT 17.04 18.34 17.36 18.62 ;
      LAYER M2 ;
        RECT 24.94 18.34 27.52 18.62 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.18 7.4 10.46 13.6 ;
      LAYER M2 ;
        RECT 11.44 28.42 28.12 28.7 ;
      LAYER M3 ;
        RECT 10.18 13.44 10.46 28.56 ;
      LAYER M2 ;
        RECT 10.32 28.42 11.61 28.7 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 25.2 10.36 33.28 10.64 ;
      LAYER M2 ;
        RECT 12.3 28 27.26 28.28 ;
      LAYER M2 ;
        RECT 25.21 10.36 25.53 10.64 ;
      LAYER M3 ;
        RECT 25.23 10.5 25.51 28.14 ;
      LAYER M2 ;
        RECT 25.21 28 25.53 28.28 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 20.5 26.3 20.78 32.08 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 8.46 18.74 8.74 24.94 ;
      LAYER M3 ;
        RECT 28.67 8.24 28.95 14.44 ;
      LAYER M3 ;
        RECT 28.24 0.68 28.52 6.88 ;
      LAYER M3 ;
        RECT 8.46 15.54 8.74 18.9 ;
      LAYER M2 ;
        RECT 8.6 15.4 28.81 15.68 ;
      LAYER M3 ;
        RECT 28.67 14.28 28.95 15.54 ;
      LAYER M3 ;
        RECT 28.67 7.56 28.95 8.4 ;
      LAYER M2 ;
        RECT 28.38 7.42 28.81 7.7 ;
      LAYER M3 ;
        RECT 28.24 6.72 28.52 7.56 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 4.13 22.54 12.21 22.82 ;
      LAYER M2 ;
        RECT 1.12 30.1 9.2 30.38 ;
      LAYER M2 ;
        RECT 4.14 22.54 4.46 22.82 ;
      LAYER M3 ;
        RECT 4.16 22.68 4.44 30.24 ;
      LAYER M2 ;
        RECT 4.14 30.1 4.46 30.38 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 24.77 2.8 32.85 3.08 ;
      LAYER M2 ;
        RECT 17.03 22.54 25.11 22.82 ;
      LAYER M2 ;
        RECT 24.78 2.8 25.1 3.08 ;
      LAYER M3 ;
        RECT 24.8 2.94 25.08 22.68 ;
      LAYER M2 ;
        RECT 24.78 22.54 25.1 22.82 ;
    END
  END F
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 27.35 22.54 35.43 22.82 ;
      LAYER M2 ;
        RECT 30.36 30.1 38.44 30.38 ;
      LAYER M2 ;
        RECT 30.37 22.54 30.69 22.82 ;
      LAYER M3 ;
        RECT 30.39 22.68 30.67 30.24 ;
      LAYER M2 ;
        RECT 30.37 30.1 30.69 30.38 ;
    END
  END C
  OBS 
  LAYER M3 ;
        RECT 18.78 3.62 19.06 9.82 ;
  LAYER M2 ;
        RECT 24.77 7 32.85 7.28 ;
  LAYER M3 ;
        RECT 18.78 6.955 19.06 7.325 ;
  LAYER M2 ;
        RECT 18.92 7 24.94 7.28 ;
  LAYER M2 ;
        RECT 18.76 7 19.08 7.28 ;
  LAYER M3 ;
        RECT 18.78 6.98 19.06 7.3 ;
  LAYER M2 ;
        RECT 18.76 7 19.08 7.28 ;
  LAYER M3 ;
        RECT 18.78 6.98 19.06 7.3 ;
  LAYER M2 ;
        RECT 1.12 25.9 9.2 26.18 ;
  LAYER M3 ;
        RECT 21.36 18.74 21.64 24.94 ;
  LAYER M3 ;
        RECT 18.78 11.18 19.06 17.38 ;
  LAYER M2 ;
        RECT 30.36 25.9 38.44 26.18 ;
  LAYER M2 ;
        RECT 9.03 25.9 21.5 26.18 ;
  LAYER M3 ;
        RECT 21.36 24.78 21.64 26.04 ;
  LAYER M3 ;
        RECT 21.36 17.64 21.64 18.9 ;
  LAYER M2 ;
        RECT 18.92 17.5 21.5 17.78 ;
  LAYER M3 ;
        RECT 18.78 17.22 19.06 17.64 ;
  LAYER M2 ;
        RECT 21.5 25.9 30.53 26.18 ;
  LAYER M2 ;
        RECT 21.34 25.9 21.66 26.18 ;
  LAYER M3 ;
        RECT 21.36 25.88 21.64 26.2 ;
  LAYER M2 ;
        RECT 21.34 25.9 21.66 26.18 ;
  LAYER M3 ;
        RECT 21.36 25.88 21.64 26.2 ;
  LAYER M2 ;
        RECT 18.76 17.5 19.08 17.78 ;
  LAYER M3 ;
        RECT 18.78 17.48 19.06 17.8 ;
  LAYER M2 ;
        RECT 21.34 17.5 21.66 17.78 ;
  LAYER M3 ;
        RECT 21.36 17.48 21.64 17.8 ;
  LAYER M2 ;
        RECT 21.34 25.9 21.66 26.18 ;
  LAYER M3 ;
        RECT 21.36 25.88 21.64 26.2 ;
  LAYER M2 ;
        RECT 18.76 17.5 19.08 17.78 ;
  LAYER M3 ;
        RECT 18.78 17.48 19.06 17.8 ;
  LAYER M2 ;
        RECT 21.34 17.5 21.66 17.78 ;
  LAYER M3 ;
        RECT 21.36 17.48 21.64 17.8 ;
  LAYER M2 ;
        RECT 21.34 25.9 21.66 26.18 ;
  LAYER M3 ;
        RECT 21.36 25.88 21.64 26.2 ;
  LAYER M2 ;
        RECT 18.76 17.5 19.08 17.78 ;
  LAYER M3 ;
        RECT 18.78 17.48 19.06 17.8 ;
  LAYER M2 ;
        RECT 21.34 17.5 21.66 17.78 ;
  LAYER M3 ;
        RECT 21.36 17.48 21.64 17.8 ;
  LAYER M2 ;
        RECT 21.34 25.9 21.66 26.18 ;
  LAYER M3 ;
        RECT 21.36 25.88 21.64 26.2 ;
  LAYER M2 ;
        RECT 18.76 17.5 19.08 17.78 ;
  LAYER M3 ;
        RECT 18.78 17.48 19.06 17.8 ;
  LAYER M2 ;
        RECT 21.34 17.5 21.66 17.78 ;
  LAYER M3 ;
        RECT 21.36 17.48 21.64 17.8 ;
  LAYER M2 ;
        RECT 21.34 25.9 21.66 26.18 ;
  LAYER M3 ;
        RECT 21.36 25.88 21.64 26.2 ;
  LAYER M2 ;
        RECT 11.44 32.62 28.12 32.9 ;
  LAYER M3 ;
        RECT 33.83 26.3 34.11 32.5 ;
  LAYER M2 ;
        RECT 27.95 32.62 33.97 32.9 ;
  LAYER M3 ;
        RECT 33.83 32.34 34.11 32.76 ;
  LAYER M2 ;
        RECT 33.81 32.62 34.13 32.9 ;
  LAYER M3 ;
        RECT 33.83 32.6 34.11 32.92 ;
  LAYER M2 ;
        RECT 33.81 32.62 34.13 32.9 ;
  LAYER M3 ;
        RECT 33.83 32.6 34.11 32.92 ;
  LAYER M3 ;
        RECT 5.45 26.3 5.73 32.5 ;
  LAYER M2 ;
        RECT 12.3 32.2 27.26 32.48 ;
  LAYER M3 ;
        RECT 5.45 31.735 5.73 32.105 ;
  LAYER M2 ;
        RECT 5.59 31.78 10.32 32.06 ;
  LAYER M1 ;
        RECT 10.195 31.92 10.445 32.34 ;
  LAYER M2 ;
        RECT 10.32 32.2 12.47 32.48 ;
  LAYER M1 ;
        RECT 10.195 31.835 10.445 32.005 ;
  LAYER M2 ;
        RECT 10.15 31.78 10.49 32.06 ;
  LAYER M1 ;
        RECT 10.195 32.255 10.445 32.425 ;
  LAYER M2 ;
        RECT 10.15 32.2 10.49 32.48 ;
  LAYER M2 ;
        RECT 5.43 31.78 5.75 32.06 ;
  LAYER M3 ;
        RECT 5.45 31.76 5.73 32.08 ;
  LAYER M1 ;
        RECT 10.195 31.835 10.445 32.005 ;
  LAYER M2 ;
        RECT 10.15 31.78 10.49 32.06 ;
  LAYER M1 ;
        RECT 10.195 32.255 10.445 32.425 ;
  LAYER M2 ;
        RECT 10.15 32.2 10.49 32.48 ;
  LAYER M2 ;
        RECT 5.43 31.78 5.75 32.06 ;
  LAYER M3 ;
        RECT 5.45 31.76 5.73 32.08 ;
  LAYER M3 ;
        RECT 10.61 5.3 10.89 17.38 ;
  LAYER M2 ;
        RECT 4.13 18.34 12.21 18.62 ;
  LAYER M2 ;
        RECT 25.2 14.56 33.28 14.84 ;
  LAYER M3 ;
        RECT 30.82 18.74 31.1 24.94 ;
  LAYER M3 ;
        RECT 10.61 17.22 10.89 18.48 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 14.515 10.89 14.885 ;
  LAYER M2 ;
        RECT 10.75 14.56 25.37 14.84 ;
  LAYER M2 ;
        RECT 30.8 14.56 31.12 14.84 ;
  LAYER M3 ;
        RECT 30.82 14.7 31.1 18.9 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 18.32 10.89 18.64 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 18.32 10.89 18.64 ;
  LAYER M2 ;
        RECT 10.59 14.56 10.91 14.84 ;
  LAYER M3 ;
        RECT 10.61 14.54 10.89 14.86 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 18.32 10.89 18.64 ;
  LAYER M2 ;
        RECT 10.59 14.56 10.91 14.84 ;
  LAYER M3 ;
        RECT 10.61 14.54 10.89 14.86 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 18.32 10.89 18.64 ;
  LAYER M2 ;
        RECT 10.59 14.56 10.91 14.84 ;
  LAYER M3 ;
        RECT 10.61 14.54 10.89 14.86 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 18.32 10.89 18.64 ;
  LAYER M2 ;
        RECT 30.8 14.56 31.12 14.84 ;
  LAYER M3 ;
        RECT 30.82 14.54 31.1 14.86 ;
  LAYER M2 ;
        RECT 10.59 14.56 10.91 14.84 ;
  LAYER M3 ;
        RECT 10.61 14.54 10.89 14.86 ;
  LAYER M2 ;
        RECT 10.59 18.34 10.91 18.62 ;
  LAYER M3 ;
        RECT 10.61 18.32 10.89 18.64 ;
  LAYER M2 ;
        RECT 30.8 14.56 31.12 14.84 ;
  LAYER M3 ;
        RECT 30.82 14.54 31.1 14.86 ;
  LAYER M1 ;
        RECT 14.495 6.635 14.745 10.165 ;
  LAYER M1 ;
        RECT 14.495 5.375 14.745 6.385 ;
  LAYER M1 ;
        RECT 14.495 3.275 14.745 4.285 ;
  LAYER M1 ;
        RECT 14.065 6.635 14.315 10.165 ;
  LAYER M1 ;
        RECT 14.925 6.635 15.175 10.165 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 10.165 ;
  LAYER M1 ;
        RECT 15.355 5.375 15.605 6.385 ;
  LAYER M1 ;
        RECT 15.355 3.275 15.605 4.285 ;
  LAYER M1 ;
        RECT 15.785 6.635 16.035 10.165 ;
  LAYER M1 ;
        RECT 16.215 6.635 16.465 10.165 ;
  LAYER M1 ;
        RECT 16.215 5.375 16.465 6.385 ;
  LAYER M1 ;
        RECT 16.215 3.275 16.465 4.285 ;
  LAYER M1 ;
        RECT 16.645 6.635 16.895 10.165 ;
  LAYER M1 ;
        RECT 17.075 6.635 17.325 10.165 ;
  LAYER M1 ;
        RECT 17.075 5.375 17.325 6.385 ;
  LAYER M1 ;
        RECT 17.075 3.275 17.325 4.285 ;
  LAYER M1 ;
        RECT 17.505 6.635 17.755 10.165 ;
  LAYER M1 ;
        RECT 17.935 6.635 18.185 10.165 ;
  LAYER M1 ;
        RECT 17.935 5.375 18.185 6.385 ;
  LAYER M1 ;
        RECT 17.935 3.275 18.185 4.285 ;
  LAYER M1 ;
        RECT 18.365 6.635 18.615 10.165 ;
  LAYER M1 ;
        RECT 18.795 6.635 19.045 10.165 ;
  LAYER M1 ;
        RECT 18.795 5.375 19.045 6.385 ;
  LAYER M1 ;
        RECT 18.795 3.275 19.045 4.285 ;
  LAYER M1 ;
        RECT 19.225 6.635 19.475 10.165 ;
  LAYER M1 ;
        RECT 19.655 6.635 19.905 10.165 ;
  LAYER M1 ;
        RECT 19.655 5.375 19.905 6.385 ;
  LAYER M1 ;
        RECT 19.655 3.275 19.905 4.285 ;
  LAYER M1 ;
        RECT 20.085 6.635 20.335 10.165 ;
  LAYER M1 ;
        RECT 20.515 6.635 20.765 10.165 ;
  LAYER M1 ;
        RECT 20.515 5.375 20.765 6.385 ;
  LAYER M1 ;
        RECT 20.515 3.275 20.765 4.285 ;
  LAYER M1 ;
        RECT 20.945 6.635 21.195 10.165 ;
  LAYER M1 ;
        RECT 21.375 6.635 21.625 10.165 ;
  LAYER M1 ;
        RECT 21.375 5.375 21.625 6.385 ;
  LAYER M1 ;
        RECT 21.375 3.275 21.625 4.285 ;
  LAYER M1 ;
        RECT 21.805 6.635 22.055 10.165 ;
  LAYER M1 ;
        RECT 22.235 6.635 22.485 10.165 ;
  LAYER M1 ;
        RECT 22.235 5.375 22.485 6.385 ;
  LAYER M1 ;
        RECT 22.235 3.275 22.485 4.285 ;
  LAYER M1 ;
        RECT 22.665 6.635 22.915 10.165 ;
  LAYER M2 ;
        RECT 14.45 3.64 22.53 3.92 ;
  LAYER M2 ;
        RECT 14.02 9.52 22.96 9.8 ;
  LAYER M2 ;
        RECT 14.45 9.94 22.53 10.22 ;
  LAYER M2 ;
        RECT 14.45 5.74 22.53 6.02 ;
  LAYER M3 ;
        RECT 18.78 3.62 19.06 9.82 ;
  LAYER M1 ;
        RECT 14.495 10.835 14.745 14.365 ;
  LAYER M1 ;
        RECT 14.495 14.615 14.745 15.625 ;
  LAYER M1 ;
        RECT 14.495 16.715 14.745 17.725 ;
  LAYER M1 ;
        RECT 14.065 10.835 14.315 14.365 ;
  LAYER M1 ;
        RECT 14.925 10.835 15.175 14.365 ;
  LAYER M1 ;
        RECT 15.355 10.835 15.605 14.365 ;
  LAYER M1 ;
        RECT 15.355 14.615 15.605 15.625 ;
  LAYER M1 ;
        RECT 15.355 16.715 15.605 17.725 ;
  LAYER M1 ;
        RECT 15.785 10.835 16.035 14.365 ;
  LAYER M1 ;
        RECT 16.215 10.835 16.465 14.365 ;
  LAYER M1 ;
        RECT 16.215 14.615 16.465 15.625 ;
  LAYER M1 ;
        RECT 16.215 16.715 16.465 17.725 ;
  LAYER M1 ;
        RECT 16.645 10.835 16.895 14.365 ;
  LAYER M1 ;
        RECT 17.075 10.835 17.325 14.365 ;
  LAYER M1 ;
        RECT 17.075 14.615 17.325 15.625 ;
  LAYER M1 ;
        RECT 17.075 16.715 17.325 17.725 ;
  LAYER M1 ;
        RECT 17.505 10.835 17.755 14.365 ;
  LAYER M1 ;
        RECT 17.935 10.835 18.185 14.365 ;
  LAYER M1 ;
        RECT 17.935 14.615 18.185 15.625 ;
  LAYER M1 ;
        RECT 17.935 16.715 18.185 17.725 ;
  LAYER M1 ;
        RECT 18.365 10.835 18.615 14.365 ;
  LAYER M1 ;
        RECT 18.795 10.835 19.045 14.365 ;
  LAYER M1 ;
        RECT 18.795 14.615 19.045 15.625 ;
  LAYER M1 ;
        RECT 18.795 16.715 19.045 17.725 ;
  LAYER M1 ;
        RECT 19.225 10.835 19.475 14.365 ;
  LAYER M1 ;
        RECT 19.655 10.835 19.905 14.365 ;
  LAYER M1 ;
        RECT 19.655 14.615 19.905 15.625 ;
  LAYER M1 ;
        RECT 19.655 16.715 19.905 17.725 ;
  LAYER M1 ;
        RECT 20.085 10.835 20.335 14.365 ;
  LAYER M1 ;
        RECT 20.515 10.835 20.765 14.365 ;
  LAYER M1 ;
        RECT 20.515 14.615 20.765 15.625 ;
  LAYER M1 ;
        RECT 20.515 16.715 20.765 17.725 ;
  LAYER M1 ;
        RECT 20.945 10.835 21.195 14.365 ;
  LAYER M1 ;
        RECT 21.375 10.835 21.625 14.365 ;
  LAYER M1 ;
        RECT 21.375 14.615 21.625 15.625 ;
  LAYER M1 ;
        RECT 21.375 16.715 21.625 17.725 ;
  LAYER M1 ;
        RECT 21.805 10.835 22.055 14.365 ;
  LAYER M1 ;
        RECT 22.235 10.835 22.485 14.365 ;
  LAYER M1 ;
        RECT 22.235 14.615 22.485 15.625 ;
  LAYER M1 ;
        RECT 22.235 16.715 22.485 17.725 ;
  LAYER M1 ;
        RECT 22.665 10.835 22.915 14.365 ;
  LAYER M2 ;
        RECT 14.45 17.08 22.53 17.36 ;
  LAYER M2 ;
        RECT 14.02 11.2 22.96 11.48 ;
  LAYER M2 ;
        RECT 14.45 10.78 22.53 11.06 ;
  LAYER M2 ;
        RECT 14.45 14.98 22.53 15.26 ;
  LAYER M3 ;
        RECT 18.78 11.18 19.06 17.38 ;
  LAYER M1 ;
        RECT 11.485 29.315 11.735 32.845 ;
  LAYER M1 ;
        RECT 11.485 28.055 11.735 29.065 ;
  LAYER M1 ;
        RECT 11.485 25.955 11.735 26.965 ;
  LAYER M1 ;
        RECT 11.055 29.315 11.305 32.845 ;
  LAYER M1 ;
        RECT 11.915 29.315 12.165 32.845 ;
  LAYER M1 ;
        RECT 12.345 29.315 12.595 32.845 ;
  LAYER M1 ;
        RECT 12.345 28.055 12.595 29.065 ;
  LAYER M1 ;
        RECT 12.345 25.955 12.595 26.965 ;
  LAYER M1 ;
        RECT 12.775 29.315 13.025 32.845 ;
  LAYER M1 ;
        RECT 13.205 29.315 13.455 32.845 ;
  LAYER M1 ;
        RECT 13.205 28.055 13.455 29.065 ;
  LAYER M1 ;
        RECT 13.205 25.955 13.455 26.965 ;
  LAYER M1 ;
        RECT 13.635 29.315 13.885 32.845 ;
  LAYER M1 ;
        RECT 14.065 29.315 14.315 32.845 ;
  LAYER M1 ;
        RECT 14.065 28.055 14.315 29.065 ;
  LAYER M1 ;
        RECT 14.065 25.955 14.315 26.965 ;
  LAYER M1 ;
        RECT 14.495 29.315 14.745 32.845 ;
  LAYER M1 ;
        RECT 14.925 29.315 15.175 32.845 ;
  LAYER M1 ;
        RECT 14.925 28.055 15.175 29.065 ;
  LAYER M1 ;
        RECT 14.925 25.955 15.175 26.965 ;
  LAYER M1 ;
        RECT 15.355 29.315 15.605 32.845 ;
  LAYER M1 ;
        RECT 15.785 29.315 16.035 32.845 ;
  LAYER M1 ;
        RECT 15.785 28.055 16.035 29.065 ;
  LAYER M1 ;
        RECT 15.785 25.955 16.035 26.965 ;
  LAYER M1 ;
        RECT 16.215 29.315 16.465 32.845 ;
  LAYER M1 ;
        RECT 16.645 29.315 16.895 32.845 ;
  LAYER M1 ;
        RECT 16.645 28.055 16.895 29.065 ;
  LAYER M1 ;
        RECT 16.645 25.955 16.895 26.965 ;
  LAYER M1 ;
        RECT 17.075 29.315 17.325 32.845 ;
  LAYER M1 ;
        RECT 17.505 29.315 17.755 32.845 ;
  LAYER M1 ;
        RECT 17.505 28.055 17.755 29.065 ;
  LAYER M1 ;
        RECT 17.505 25.955 17.755 26.965 ;
  LAYER M1 ;
        RECT 17.935 29.315 18.185 32.845 ;
  LAYER M1 ;
        RECT 18.365 29.315 18.615 32.845 ;
  LAYER M1 ;
        RECT 18.365 28.055 18.615 29.065 ;
  LAYER M1 ;
        RECT 18.365 25.955 18.615 26.965 ;
  LAYER M1 ;
        RECT 18.795 29.315 19.045 32.845 ;
  LAYER M1 ;
        RECT 19.225 29.315 19.475 32.845 ;
  LAYER M1 ;
        RECT 19.225 28.055 19.475 29.065 ;
  LAYER M1 ;
        RECT 19.225 25.955 19.475 26.965 ;
  LAYER M1 ;
        RECT 19.655 29.315 19.905 32.845 ;
  LAYER M1 ;
        RECT 20.085 29.315 20.335 32.845 ;
  LAYER M1 ;
        RECT 20.085 28.055 20.335 29.065 ;
  LAYER M1 ;
        RECT 20.085 25.955 20.335 26.965 ;
  LAYER M1 ;
        RECT 20.515 29.315 20.765 32.845 ;
  LAYER M1 ;
        RECT 20.945 29.315 21.195 32.845 ;
  LAYER M1 ;
        RECT 20.945 28.055 21.195 29.065 ;
  LAYER M1 ;
        RECT 20.945 25.955 21.195 26.965 ;
  LAYER M1 ;
        RECT 21.375 29.315 21.625 32.845 ;
  LAYER M1 ;
        RECT 21.805 29.315 22.055 32.845 ;
  LAYER M1 ;
        RECT 21.805 28.055 22.055 29.065 ;
  LAYER M1 ;
        RECT 21.805 25.955 22.055 26.965 ;
  LAYER M1 ;
        RECT 22.235 29.315 22.485 32.845 ;
  LAYER M1 ;
        RECT 22.665 29.315 22.915 32.845 ;
  LAYER M1 ;
        RECT 22.665 28.055 22.915 29.065 ;
  LAYER M1 ;
        RECT 22.665 25.955 22.915 26.965 ;
  LAYER M1 ;
        RECT 23.095 29.315 23.345 32.845 ;
  LAYER M1 ;
        RECT 23.525 29.315 23.775 32.845 ;
  LAYER M1 ;
        RECT 23.525 28.055 23.775 29.065 ;
  LAYER M1 ;
        RECT 23.525 25.955 23.775 26.965 ;
  LAYER M1 ;
        RECT 23.955 29.315 24.205 32.845 ;
  LAYER M1 ;
        RECT 24.385 29.315 24.635 32.845 ;
  LAYER M1 ;
        RECT 24.385 28.055 24.635 29.065 ;
  LAYER M1 ;
        RECT 24.385 25.955 24.635 26.965 ;
  LAYER M1 ;
        RECT 24.815 29.315 25.065 32.845 ;
  LAYER M1 ;
        RECT 25.245 29.315 25.495 32.845 ;
  LAYER M1 ;
        RECT 25.245 28.055 25.495 29.065 ;
  LAYER M1 ;
        RECT 25.245 25.955 25.495 26.965 ;
  LAYER M1 ;
        RECT 25.675 29.315 25.925 32.845 ;
  LAYER M1 ;
        RECT 26.105 29.315 26.355 32.845 ;
  LAYER M1 ;
        RECT 26.105 28.055 26.355 29.065 ;
  LAYER M1 ;
        RECT 26.105 25.955 26.355 26.965 ;
  LAYER M1 ;
        RECT 26.535 29.315 26.785 32.845 ;
  LAYER M1 ;
        RECT 26.965 29.315 27.215 32.845 ;
  LAYER M1 ;
        RECT 26.965 28.055 27.215 29.065 ;
  LAYER M1 ;
        RECT 26.965 25.955 27.215 26.965 ;
  LAYER M1 ;
        RECT 27.395 29.315 27.645 32.845 ;
  LAYER M1 ;
        RECT 27.825 29.315 28.075 32.845 ;
  LAYER M1 ;
        RECT 27.825 28.055 28.075 29.065 ;
  LAYER M1 ;
        RECT 27.825 25.955 28.075 26.965 ;
  LAYER M1 ;
        RECT 28.255 29.315 28.505 32.845 ;
  LAYER M2 ;
        RECT 11.44 26.32 28.12 26.6 ;
  LAYER M2 ;
        RECT 11.01 31.78 28.55 32.06 ;
  LAYER M2 ;
        RECT 11.44 32.62 28.12 32.9 ;
  LAYER M2 ;
        RECT 12.3 32.2 27.26 32.48 ;
  LAYER M2 ;
        RECT 11.44 28.42 28.12 28.7 ;
  LAYER M2 ;
        RECT 12.3 28 27.26 28.28 ;
  LAYER M3 ;
        RECT 20.5 26.3 20.78 32.08 ;
  LAYER M1 ;
        RECT 32.985 11.255 33.235 14.785 ;
  LAYER M1 ;
        RECT 32.985 9.995 33.235 11.005 ;
  LAYER M1 ;
        RECT 32.985 7.895 33.235 8.905 ;
  LAYER M1 ;
        RECT 33.415 11.255 33.665 14.785 ;
  LAYER M1 ;
        RECT 32.555 11.255 32.805 14.785 ;
  LAYER M1 ;
        RECT 32.125 11.255 32.375 14.785 ;
  LAYER M1 ;
        RECT 32.125 9.995 32.375 11.005 ;
  LAYER M1 ;
        RECT 32.125 7.895 32.375 8.905 ;
  LAYER M1 ;
        RECT 31.695 11.255 31.945 14.785 ;
  LAYER M1 ;
        RECT 31.265 11.255 31.515 14.785 ;
  LAYER M1 ;
        RECT 31.265 9.995 31.515 11.005 ;
  LAYER M1 ;
        RECT 31.265 7.895 31.515 8.905 ;
  LAYER M1 ;
        RECT 30.835 11.255 31.085 14.785 ;
  LAYER M1 ;
        RECT 30.405 11.255 30.655 14.785 ;
  LAYER M1 ;
        RECT 30.405 9.995 30.655 11.005 ;
  LAYER M1 ;
        RECT 30.405 7.895 30.655 8.905 ;
  LAYER M1 ;
        RECT 29.975 11.255 30.225 14.785 ;
  LAYER M1 ;
        RECT 29.545 11.255 29.795 14.785 ;
  LAYER M1 ;
        RECT 29.545 9.995 29.795 11.005 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 8.905 ;
  LAYER M1 ;
        RECT 29.115 11.255 29.365 14.785 ;
  LAYER M1 ;
        RECT 28.685 11.255 28.935 14.785 ;
  LAYER M1 ;
        RECT 28.685 9.995 28.935 11.005 ;
  LAYER M1 ;
        RECT 28.685 7.895 28.935 8.905 ;
  LAYER M1 ;
        RECT 28.255 11.255 28.505 14.785 ;
  LAYER M1 ;
        RECT 27.825 11.255 28.075 14.785 ;
  LAYER M1 ;
        RECT 27.825 9.995 28.075 11.005 ;
  LAYER M1 ;
        RECT 27.825 7.895 28.075 8.905 ;
  LAYER M1 ;
        RECT 27.395 11.255 27.645 14.785 ;
  LAYER M1 ;
        RECT 26.965 11.255 27.215 14.785 ;
  LAYER M1 ;
        RECT 26.965 9.995 27.215 11.005 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 8.905 ;
  LAYER M1 ;
        RECT 26.535 11.255 26.785 14.785 ;
  LAYER M1 ;
        RECT 26.105 11.255 26.355 14.785 ;
  LAYER M1 ;
        RECT 26.105 9.995 26.355 11.005 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 8.905 ;
  LAYER M1 ;
        RECT 25.675 11.255 25.925 14.785 ;
  LAYER M1 ;
        RECT 25.245 11.255 25.495 14.785 ;
  LAYER M1 ;
        RECT 25.245 9.995 25.495 11.005 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 8.905 ;
  LAYER M1 ;
        RECT 24.815 11.255 25.065 14.785 ;
  LAYER M2 ;
        RECT 25.2 8.26 33.28 8.54 ;
  LAYER M2 ;
        RECT 24.77 14.14 33.71 14.42 ;
  LAYER M2 ;
        RECT 25.2 14.56 33.28 14.84 ;
  LAYER M2 ;
        RECT 25.2 10.36 33.28 10.64 ;
  LAYER M3 ;
        RECT 28.67 8.24 28.95 14.44 ;
  LAYER M1 ;
        RECT 4.175 18.395 4.425 21.925 ;
  LAYER M1 ;
        RECT 4.175 22.175 4.425 23.185 ;
  LAYER M1 ;
        RECT 4.175 24.275 4.425 25.285 ;
  LAYER M1 ;
        RECT 3.745 18.395 3.995 21.925 ;
  LAYER M1 ;
        RECT 4.605 18.395 4.855 21.925 ;
  LAYER M1 ;
        RECT 5.035 18.395 5.285 21.925 ;
  LAYER M1 ;
        RECT 5.035 22.175 5.285 23.185 ;
  LAYER M1 ;
        RECT 5.035 24.275 5.285 25.285 ;
  LAYER M1 ;
        RECT 5.465 18.395 5.715 21.925 ;
  LAYER M1 ;
        RECT 5.895 18.395 6.145 21.925 ;
  LAYER M1 ;
        RECT 5.895 22.175 6.145 23.185 ;
  LAYER M1 ;
        RECT 5.895 24.275 6.145 25.285 ;
  LAYER M1 ;
        RECT 6.325 18.395 6.575 21.925 ;
  LAYER M1 ;
        RECT 6.755 18.395 7.005 21.925 ;
  LAYER M1 ;
        RECT 6.755 22.175 7.005 23.185 ;
  LAYER M1 ;
        RECT 6.755 24.275 7.005 25.285 ;
  LAYER M1 ;
        RECT 7.185 18.395 7.435 21.925 ;
  LAYER M1 ;
        RECT 7.615 18.395 7.865 21.925 ;
  LAYER M1 ;
        RECT 7.615 22.175 7.865 23.185 ;
  LAYER M1 ;
        RECT 7.615 24.275 7.865 25.285 ;
  LAYER M1 ;
        RECT 8.045 18.395 8.295 21.925 ;
  LAYER M1 ;
        RECT 8.475 18.395 8.725 21.925 ;
  LAYER M1 ;
        RECT 8.475 22.175 8.725 23.185 ;
  LAYER M1 ;
        RECT 8.475 24.275 8.725 25.285 ;
  LAYER M1 ;
        RECT 8.905 18.395 9.155 21.925 ;
  LAYER M1 ;
        RECT 9.335 18.395 9.585 21.925 ;
  LAYER M1 ;
        RECT 9.335 22.175 9.585 23.185 ;
  LAYER M1 ;
        RECT 9.335 24.275 9.585 25.285 ;
  LAYER M1 ;
        RECT 9.765 18.395 10.015 21.925 ;
  LAYER M1 ;
        RECT 10.195 18.395 10.445 21.925 ;
  LAYER M1 ;
        RECT 10.195 22.175 10.445 23.185 ;
  LAYER M1 ;
        RECT 10.195 24.275 10.445 25.285 ;
  LAYER M1 ;
        RECT 10.625 18.395 10.875 21.925 ;
  LAYER M1 ;
        RECT 11.055 18.395 11.305 21.925 ;
  LAYER M1 ;
        RECT 11.055 22.175 11.305 23.185 ;
  LAYER M1 ;
        RECT 11.055 24.275 11.305 25.285 ;
  LAYER M1 ;
        RECT 11.485 18.395 11.735 21.925 ;
  LAYER M1 ;
        RECT 11.915 18.395 12.165 21.925 ;
  LAYER M1 ;
        RECT 11.915 22.175 12.165 23.185 ;
  LAYER M1 ;
        RECT 11.915 24.275 12.165 25.285 ;
  LAYER M1 ;
        RECT 12.345 18.395 12.595 21.925 ;
  LAYER M2 ;
        RECT 4.13 24.64 12.21 24.92 ;
  LAYER M2 ;
        RECT 3.7 18.76 12.64 19.04 ;
  LAYER M2 ;
        RECT 4.13 18.34 12.21 18.62 ;
  LAYER M2 ;
        RECT 4.13 22.54 12.21 22.82 ;
  LAYER M3 ;
        RECT 8.46 18.74 8.74 24.94 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.555 2.435 32.805 3.445 ;
  LAYER M1 ;
        RECT 32.555 0.335 32.805 1.345 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 31.695 2.435 31.945 3.445 ;
  LAYER M1 ;
        RECT 31.695 0.335 31.945 1.345 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 30.835 2.435 31.085 3.445 ;
  LAYER M1 ;
        RECT 30.835 0.335 31.085 1.345 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 29.975 2.435 30.225 3.445 ;
  LAYER M1 ;
        RECT 29.975 0.335 30.225 1.345 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.115 2.435 29.365 3.445 ;
  LAYER M1 ;
        RECT 29.115 0.335 29.365 1.345 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 28.255 2.435 28.505 3.445 ;
  LAYER M1 ;
        RECT 28.255 0.335 28.505 1.345 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 27.395 2.435 27.645 3.445 ;
  LAYER M1 ;
        RECT 27.395 0.335 27.645 1.345 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.535 2.435 26.785 3.445 ;
  LAYER M1 ;
        RECT 26.535 0.335 26.785 1.345 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 25.675 2.435 25.925 3.445 ;
  LAYER M1 ;
        RECT 25.675 0.335 25.925 1.345 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 24.815 2.435 25.065 3.445 ;
  LAYER M1 ;
        RECT 24.815 0.335 25.065 1.345 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M2 ;
        RECT 24.77 0.7 32.85 0.98 ;
  LAYER M2 ;
        RECT 24.34 6.58 33.28 6.86 ;
  LAYER M2 ;
        RECT 24.77 7 32.85 7.28 ;
  LAYER M2 ;
        RECT 24.77 2.8 32.85 3.08 ;
  LAYER M3 ;
        RECT 28.24 0.68 28.52 6.88 ;
  LAYER M1 ;
        RECT 8.475 14.195 8.725 17.725 ;
  LAYER M1 ;
        RECT 8.475 12.935 8.725 13.945 ;
  LAYER M1 ;
        RECT 8.475 8.315 8.725 11.845 ;
  LAYER M1 ;
        RECT 8.475 7.055 8.725 8.065 ;
  LAYER M1 ;
        RECT 8.475 4.955 8.725 5.965 ;
  LAYER M1 ;
        RECT 8.045 14.195 8.295 17.725 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 11.845 ;
  LAYER M1 ;
        RECT 8.905 14.195 9.155 17.725 ;
  LAYER M1 ;
        RECT 8.905 8.315 9.155 11.845 ;
  LAYER M1 ;
        RECT 9.335 14.195 9.585 17.725 ;
  LAYER M1 ;
        RECT 9.335 12.935 9.585 13.945 ;
  LAYER M1 ;
        RECT 9.335 8.315 9.585 11.845 ;
  LAYER M1 ;
        RECT 9.335 7.055 9.585 8.065 ;
  LAYER M1 ;
        RECT 9.335 4.955 9.585 5.965 ;
  LAYER M1 ;
        RECT 9.765 14.195 10.015 17.725 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 11.845 ;
  LAYER M1 ;
        RECT 10.195 14.195 10.445 17.725 ;
  LAYER M1 ;
        RECT 10.195 12.935 10.445 13.945 ;
  LAYER M1 ;
        RECT 10.195 8.315 10.445 11.845 ;
  LAYER M1 ;
        RECT 10.195 7.055 10.445 8.065 ;
  LAYER M1 ;
        RECT 10.195 4.955 10.445 5.965 ;
  LAYER M1 ;
        RECT 10.625 14.195 10.875 17.725 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 11.845 ;
  LAYER M1 ;
        RECT 11.055 14.195 11.305 17.725 ;
  LAYER M1 ;
        RECT 11.055 12.935 11.305 13.945 ;
  LAYER M1 ;
        RECT 11.055 8.315 11.305 11.845 ;
  LAYER M1 ;
        RECT 11.055 7.055 11.305 8.065 ;
  LAYER M1 ;
        RECT 11.055 4.955 11.305 5.965 ;
  LAYER M1 ;
        RECT 11.485 14.195 11.735 17.725 ;
  LAYER M1 ;
        RECT 11.485 8.315 11.735 11.845 ;
  LAYER M1 ;
        RECT 11.915 14.195 12.165 17.725 ;
  LAYER M1 ;
        RECT 11.915 12.935 12.165 13.945 ;
  LAYER M1 ;
        RECT 11.915 8.315 12.165 11.845 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 8.065 ;
  LAYER M1 ;
        RECT 11.915 4.955 12.165 5.965 ;
  LAYER M1 ;
        RECT 12.345 14.195 12.595 17.725 ;
  LAYER M1 ;
        RECT 12.345 8.315 12.595 11.845 ;
  LAYER M2 ;
        RECT 8.43 17.5 12.21 17.78 ;
  LAYER M2 ;
        RECT 8.43 13.3 12.21 13.58 ;
  LAYER M2 ;
        RECT 8 17.08 12.64 17.36 ;
  LAYER M2 ;
        RECT 8.43 11.62 12.21 11.9 ;
  LAYER M2 ;
        RECT 8.43 7.42 12.21 7.7 ;
  LAYER M2 ;
        RECT 8.43 5.32 12.21 5.6 ;
  LAYER M2 ;
        RECT 8 11.2 12.64 11.48 ;
  LAYER M3 ;
        RECT 9.75 11.6 10.03 17.8 ;
  LAYER M3 ;
        RECT 10.18 7.4 10.46 13.6 ;
  LAYER M3 ;
        RECT 10.61 5.3 10.89 17.38 ;
  LAYER M1 ;
        RECT 35.135 18.395 35.385 21.925 ;
  LAYER M1 ;
        RECT 35.135 22.175 35.385 23.185 ;
  LAYER M1 ;
        RECT 35.135 24.275 35.385 25.285 ;
  LAYER M1 ;
        RECT 35.565 18.395 35.815 21.925 ;
  LAYER M1 ;
        RECT 34.705 18.395 34.955 21.925 ;
  LAYER M1 ;
        RECT 34.275 18.395 34.525 21.925 ;
  LAYER M1 ;
        RECT 34.275 22.175 34.525 23.185 ;
  LAYER M1 ;
        RECT 34.275 24.275 34.525 25.285 ;
  LAYER M1 ;
        RECT 33.845 18.395 34.095 21.925 ;
  LAYER M1 ;
        RECT 33.415 18.395 33.665 21.925 ;
  LAYER M1 ;
        RECT 33.415 22.175 33.665 23.185 ;
  LAYER M1 ;
        RECT 33.415 24.275 33.665 25.285 ;
  LAYER M1 ;
        RECT 32.985 18.395 33.235 21.925 ;
  LAYER M1 ;
        RECT 32.555 18.395 32.805 21.925 ;
  LAYER M1 ;
        RECT 32.555 22.175 32.805 23.185 ;
  LAYER M1 ;
        RECT 32.555 24.275 32.805 25.285 ;
  LAYER M1 ;
        RECT 32.125 18.395 32.375 21.925 ;
  LAYER M1 ;
        RECT 31.695 18.395 31.945 21.925 ;
  LAYER M1 ;
        RECT 31.695 22.175 31.945 23.185 ;
  LAYER M1 ;
        RECT 31.695 24.275 31.945 25.285 ;
  LAYER M1 ;
        RECT 31.265 18.395 31.515 21.925 ;
  LAYER M1 ;
        RECT 30.835 18.395 31.085 21.925 ;
  LAYER M1 ;
        RECT 30.835 22.175 31.085 23.185 ;
  LAYER M1 ;
        RECT 30.835 24.275 31.085 25.285 ;
  LAYER M1 ;
        RECT 30.405 18.395 30.655 21.925 ;
  LAYER M1 ;
        RECT 29.975 18.395 30.225 21.925 ;
  LAYER M1 ;
        RECT 29.975 22.175 30.225 23.185 ;
  LAYER M1 ;
        RECT 29.975 24.275 30.225 25.285 ;
  LAYER M1 ;
        RECT 29.545 18.395 29.795 21.925 ;
  LAYER M1 ;
        RECT 29.115 18.395 29.365 21.925 ;
  LAYER M1 ;
        RECT 29.115 22.175 29.365 23.185 ;
  LAYER M1 ;
        RECT 29.115 24.275 29.365 25.285 ;
  LAYER M1 ;
        RECT 28.685 18.395 28.935 21.925 ;
  LAYER M1 ;
        RECT 28.255 18.395 28.505 21.925 ;
  LAYER M1 ;
        RECT 28.255 22.175 28.505 23.185 ;
  LAYER M1 ;
        RECT 28.255 24.275 28.505 25.285 ;
  LAYER M1 ;
        RECT 27.825 18.395 28.075 21.925 ;
  LAYER M1 ;
        RECT 27.395 18.395 27.645 21.925 ;
  LAYER M1 ;
        RECT 27.395 22.175 27.645 23.185 ;
  LAYER M1 ;
        RECT 27.395 24.275 27.645 25.285 ;
  LAYER M1 ;
        RECT 26.965 18.395 27.215 21.925 ;
  LAYER M2 ;
        RECT 27.35 24.64 35.43 24.92 ;
  LAYER M2 ;
        RECT 26.92 18.76 35.86 19.04 ;
  LAYER M2 ;
        RECT 27.35 18.34 35.43 18.62 ;
  LAYER M2 ;
        RECT 27.35 22.54 35.43 22.82 ;
  LAYER M3 ;
        RECT 30.82 18.74 31.1 24.94 ;
  LAYER M1 ;
        RECT 38.145 25.955 38.395 29.485 ;
  LAYER M1 ;
        RECT 38.145 29.735 38.395 30.745 ;
  LAYER M1 ;
        RECT 38.145 31.835 38.395 32.845 ;
  LAYER M1 ;
        RECT 38.575 25.955 38.825 29.485 ;
  LAYER M1 ;
        RECT 37.715 25.955 37.965 29.485 ;
  LAYER M1 ;
        RECT 37.285 25.955 37.535 29.485 ;
  LAYER M1 ;
        RECT 37.285 29.735 37.535 30.745 ;
  LAYER M1 ;
        RECT 37.285 31.835 37.535 32.845 ;
  LAYER M1 ;
        RECT 36.855 25.955 37.105 29.485 ;
  LAYER M1 ;
        RECT 36.425 25.955 36.675 29.485 ;
  LAYER M1 ;
        RECT 36.425 29.735 36.675 30.745 ;
  LAYER M1 ;
        RECT 36.425 31.835 36.675 32.845 ;
  LAYER M1 ;
        RECT 35.995 25.955 36.245 29.485 ;
  LAYER M1 ;
        RECT 35.565 25.955 35.815 29.485 ;
  LAYER M1 ;
        RECT 35.565 29.735 35.815 30.745 ;
  LAYER M1 ;
        RECT 35.565 31.835 35.815 32.845 ;
  LAYER M1 ;
        RECT 35.135 25.955 35.385 29.485 ;
  LAYER M1 ;
        RECT 34.705 25.955 34.955 29.485 ;
  LAYER M1 ;
        RECT 34.705 29.735 34.955 30.745 ;
  LAYER M1 ;
        RECT 34.705 31.835 34.955 32.845 ;
  LAYER M1 ;
        RECT 34.275 25.955 34.525 29.485 ;
  LAYER M1 ;
        RECT 33.845 25.955 34.095 29.485 ;
  LAYER M1 ;
        RECT 33.845 29.735 34.095 30.745 ;
  LAYER M1 ;
        RECT 33.845 31.835 34.095 32.845 ;
  LAYER M1 ;
        RECT 33.415 25.955 33.665 29.485 ;
  LAYER M1 ;
        RECT 32.985 25.955 33.235 29.485 ;
  LAYER M1 ;
        RECT 32.985 29.735 33.235 30.745 ;
  LAYER M1 ;
        RECT 32.985 31.835 33.235 32.845 ;
  LAYER M1 ;
        RECT 32.555 25.955 32.805 29.485 ;
  LAYER M1 ;
        RECT 32.125 25.955 32.375 29.485 ;
  LAYER M1 ;
        RECT 32.125 29.735 32.375 30.745 ;
  LAYER M1 ;
        RECT 32.125 31.835 32.375 32.845 ;
  LAYER M1 ;
        RECT 31.695 25.955 31.945 29.485 ;
  LAYER M1 ;
        RECT 31.265 25.955 31.515 29.485 ;
  LAYER M1 ;
        RECT 31.265 29.735 31.515 30.745 ;
  LAYER M1 ;
        RECT 31.265 31.835 31.515 32.845 ;
  LAYER M1 ;
        RECT 30.835 25.955 31.085 29.485 ;
  LAYER M1 ;
        RECT 30.405 25.955 30.655 29.485 ;
  LAYER M1 ;
        RECT 30.405 29.735 30.655 30.745 ;
  LAYER M1 ;
        RECT 30.405 31.835 30.655 32.845 ;
  LAYER M1 ;
        RECT 29.975 25.955 30.225 29.485 ;
  LAYER M2 ;
        RECT 30.36 32.2 38.44 32.48 ;
  LAYER M2 ;
        RECT 29.93 26.32 38.87 26.6 ;
  LAYER M2 ;
        RECT 30.36 25.9 38.44 26.18 ;
  LAYER M2 ;
        RECT 30.36 30.1 38.44 30.38 ;
  LAYER M3 ;
        RECT 33.83 26.3 34.11 32.5 ;
  LAYER M1 ;
        RECT 1.165 25.955 1.415 29.485 ;
  LAYER M1 ;
        RECT 1.165 29.735 1.415 30.745 ;
  LAYER M1 ;
        RECT 1.165 31.835 1.415 32.845 ;
  LAYER M1 ;
        RECT 0.735 25.955 0.985 29.485 ;
  LAYER M1 ;
        RECT 1.595 25.955 1.845 29.485 ;
  LAYER M1 ;
        RECT 2.025 25.955 2.275 29.485 ;
  LAYER M1 ;
        RECT 2.025 29.735 2.275 30.745 ;
  LAYER M1 ;
        RECT 2.025 31.835 2.275 32.845 ;
  LAYER M1 ;
        RECT 2.455 25.955 2.705 29.485 ;
  LAYER M1 ;
        RECT 2.885 25.955 3.135 29.485 ;
  LAYER M1 ;
        RECT 2.885 29.735 3.135 30.745 ;
  LAYER M1 ;
        RECT 2.885 31.835 3.135 32.845 ;
  LAYER M1 ;
        RECT 3.315 25.955 3.565 29.485 ;
  LAYER M1 ;
        RECT 3.745 25.955 3.995 29.485 ;
  LAYER M1 ;
        RECT 3.745 29.735 3.995 30.745 ;
  LAYER M1 ;
        RECT 3.745 31.835 3.995 32.845 ;
  LAYER M1 ;
        RECT 4.175 25.955 4.425 29.485 ;
  LAYER M1 ;
        RECT 4.605 25.955 4.855 29.485 ;
  LAYER M1 ;
        RECT 4.605 29.735 4.855 30.745 ;
  LAYER M1 ;
        RECT 4.605 31.835 4.855 32.845 ;
  LAYER M1 ;
        RECT 5.035 25.955 5.285 29.485 ;
  LAYER M1 ;
        RECT 5.465 25.955 5.715 29.485 ;
  LAYER M1 ;
        RECT 5.465 29.735 5.715 30.745 ;
  LAYER M1 ;
        RECT 5.465 31.835 5.715 32.845 ;
  LAYER M1 ;
        RECT 5.895 25.955 6.145 29.485 ;
  LAYER M1 ;
        RECT 6.325 25.955 6.575 29.485 ;
  LAYER M1 ;
        RECT 6.325 29.735 6.575 30.745 ;
  LAYER M1 ;
        RECT 6.325 31.835 6.575 32.845 ;
  LAYER M1 ;
        RECT 6.755 25.955 7.005 29.485 ;
  LAYER M1 ;
        RECT 7.185 25.955 7.435 29.485 ;
  LAYER M1 ;
        RECT 7.185 29.735 7.435 30.745 ;
  LAYER M1 ;
        RECT 7.185 31.835 7.435 32.845 ;
  LAYER M1 ;
        RECT 7.615 25.955 7.865 29.485 ;
  LAYER M1 ;
        RECT 8.045 25.955 8.295 29.485 ;
  LAYER M1 ;
        RECT 8.045 29.735 8.295 30.745 ;
  LAYER M1 ;
        RECT 8.045 31.835 8.295 32.845 ;
  LAYER M1 ;
        RECT 8.475 25.955 8.725 29.485 ;
  LAYER M1 ;
        RECT 8.905 25.955 9.155 29.485 ;
  LAYER M1 ;
        RECT 8.905 29.735 9.155 30.745 ;
  LAYER M1 ;
        RECT 8.905 31.835 9.155 32.845 ;
  LAYER M1 ;
        RECT 9.335 25.955 9.585 29.485 ;
  LAYER M2 ;
        RECT 1.12 32.2 9.2 32.48 ;
  LAYER M2 ;
        RECT 0.69 26.32 9.63 26.6 ;
  LAYER M2 ;
        RECT 1.12 25.9 9.2 26.18 ;
  LAYER M2 ;
        RECT 1.12 30.1 9.2 30.38 ;
  LAYER M3 ;
        RECT 5.45 26.3 5.73 32.5 ;
  LAYER M1 ;
        RECT 17.075 18.395 17.325 21.925 ;
  LAYER M1 ;
        RECT 17.075 22.175 17.325 23.185 ;
  LAYER M1 ;
        RECT 17.075 24.275 17.325 25.285 ;
  LAYER M1 ;
        RECT 16.645 18.395 16.895 21.925 ;
  LAYER M1 ;
        RECT 17.505 18.395 17.755 21.925 ;
  LAYER M1 ;
        RECT 17.935 18.395 18.185 21.925 ;
  LAYER M1 ;
        RECT 17.935 22.175 18.185 23.185 ;
  LAYER M1 ;
        RECT 17.935 24.275 18.185 25.285 ;
  LAYER M1 ;
        RECT 18.365 18.395 18.615 21.925 ;
  LAYER M1 ;
        RECT 18.795 18.395 19.045 21.925 ;
  LAYER M1 ;
        RECT 18.795 22.175 19.045 23.185 ;
  LAYER M1 ;
        RECT 18.795 24.275 19.045 25.285 ;
  LAYER M1 ;
        RECT 19.225 18.395 19.475 21.925 ;
  LAYER M1 ;
        RECT 19.655 18.395 19.905 21.925 ;
  LAYER M1 ;
        RECT 19.655 22.175 19.905 23.185 ;
  LAYER M1 ;
        RECT 19.655 24.275 19.905 25.285 ;
  LAYER M1 ;
        RECT 20.085 18.395 20.335 21.925 ;
  LAYER M1 ;
        RECT 20.515 18.395 20.765 21.925 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 23.185 ;
  LAYER M1 ;
        RECT 20.515 24.275 20.765 25.285 ;
  LAYER M1 ;
        RECT 20.945 18.395 21.195 21.925 ;
  LAYER M1 ;
        RECT 21.375 18.395 21.625 21.925 ;
  LAYER M1 ;
        RECT 21.375 22.175 21.625 23.185 ;
  LAYER M1 ;
        RECT 21.375 24.275 21.625 25.285 ;
  LAYER M1 ;
        RECT 21.805 18.395 22.055 21.925 ;
  LAYER M1 ;
        RECT 22.235 18.395 22.485 21.925 ;
  LAYER M1 ;
        RECT 22.235 22.175 22.485 23.185 ;
  LAYER M1 ;
        RECT 22.235 24.275 22.485 25.285 ;
  LAYER M1 ;
        RECT 22.665 18.395 22.915 21.925 ;
  LAYER M1 ;
        RECT 23.095 18.395 23.345 21.925 ;
  LAYER M1 ;
        RECT 23.095 22.175 23.345 23.185 ;
  LAYER M1 ;
        RECT 23.095 24.275 23.345 25.285 ;
  LAYER M1 ;
        RECT 23.525 18.395 23.775 21.925 ;
  LAYER M1 ;
        RECT 23.955 18.395 24.205 21.925 ;
  LAYER M1 ;
        RECT 23.955 22.175 24.205 23.185 ;
  LAYER M1 ;
        RECT 23.955 24.275 24.205 25.285 ;
  LAYER M1 ;
        RECT 24.385 18.395 24.635 21.925 ;
  LAYER M1 ;
        RECT 24.815 18.395 25.065 21.925 ;
  LAYER M1 ;
        RECT 24.815 22.175 25.065 23.185 ;
  LAYER M1 ;
        RECT 24.815 24.275 25.065 25.285 ;
  LAYER M1 ;
        RECT 25.245 18.395 25.495 21.925 ;
  LAYER M2 ;
        RECT 17.03 24.64 25.11 24.92 ;
  LAYER M2 ;
        RECT 16.6 18.76 25.54 19.04 ;
  LAYER M2 ;
        RECT 17.03 18.34 25.11 18.62 ;
  LAYER M2 ;
        RECT 17.03 22.54 25.11 22.82 ;
  LAYER M3 ;
        RECT 21.36 18.74 21.64 24.94 ;
  END 
END FN_SIM
